// de2i_150.v

// Generated using ACDS version 13.0sp1 232 at 2014.03.05.15:52:21

`timescale 1 ps / 1 ps
module de2i_150 (
		input  wire        clk_clk,              //           clk.clk
		input  wire        reset_reset_n,        //         reset.reset_n
		input  wire        switch0_export,       //       switch0.export
		output wire [7:0]  led_export,           //           led.export
		input  wire        key0_export,          //          key0.export
		input  wire        uart_rxd,             //          uart.rxd
		output wire        uart_txd,             //              .txd
		input  wire [13:0] adc_export,           //           adc.export
		output wire        cs_export,            //            cs.export
		output wire        sclk_export,          //          sclk.export
		output wire        sdin_export,          //          sdin.export
		output wire        din_export,           //           din.export
		input  wire        bclk_in_export,       //       bclk_in.export
		input  wire        lrcout_export,        //        lrcout.export
		input  wire        dout_export,          //          dout.export
		input  wire        bclk_out_export,      //      bclk_out.export
		input  wire        lrcin_export,         //         lrcin.export
		input  wire        key1_export,          //          key1.export
		input  wire        key2_export,          //          key2.export
		input  wire        key3_export,          //          key3.export
		input  wire        switch1_export,       //       switch1.export
		input  wire        switch2_export,       //       switch2.export
		input  wire        switch3_export,       //       switch3.export
		input  wire        switch4_export,       //       switch4.export
		input  wire [15:0] leftdata_export,      //      leftdata.export
		input  wire [15:0] rightdata_export,     //     rightdata.export
		input  wire        leftready_export,     //     leftready.export
		input  wire        rightready_export,    //    rightready.export
		output wire [15:0] leftsenddata_export,  //  leftsenddata.export
		output wire [15:0] rightsenddata_export, // rightsenddata.export
		output wire        clk_12mhz_c0_clk,     //  clk_12mhz_c0.clk
		input  wire        switch5_export,       //       switch5.export
		input  wire        switch6_export,       //       switch6.export
		input  wire        switch7_export,       //       switch7.export
		input  wire        switch8_export        //       switch8.export
	);

	wire         altpll_0_c0_clk;                                                                                   // altpll_0:c0 -> [adc:clk, adc_s1_translator:clk, adc_s1_translator_avalon_universal_slave_0_agent:clk, adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, bclk_in:clk, bclk_in_s1_translator:clk, bclk_in_s1_translator_avalon_universal_slave_0_agent:clk, bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, bclk_out:clk, bclk_out_s1_translator:clk, bclk_out_s1_translator_avalon_universal_slave_0_agent:clk, bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, crosser:in_clk, crosser_001:in_clk, crosser_002:out_clk, crosser_003:out_clk, cs:clk, cs_s1_translator:clk, cs_s1_translator_avalon_universal_slave_0_agent:clk, cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, din:clk, din_s1_translator:clk, din_s1_translator_avalon_universal_slave_0_agent:clk, din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dout:clk, dout_s1_translator:clk, dout_s1_translator_avalon_universal_slave_0_agent:clk, dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, id_router_020:clk, id_router_021:clk, id_router_022:clk, id_router_023:clk, id_router_024:clk, id_router_026:clk, id_router_027:clk, id_router_028:clk, id_router_029:clk, id_router_030:clk, id_router_031:clk, id_router_033:clk, id_router_034:clk, id_router_035:clk, id_router_036:clk, irq_mapper:clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, key0:clk, key0_s1_translator:clk, key0_s1_translator_avalon_universal_slave_0_agent:clk, key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, key1:clk, key1_s1_translator:clk, key1_s1_translator_avalon_universal_slave_0_agent:clk, key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, key2:clk, key2_s1_translator:clk, key2_s1_translator_avalon_universal_slave_0_agent:clk, key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, key3:clk, key3_s1_translator:clk, key3_s1_translator_avalon_universal_slave_0_agent:clk, key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, led:clk, led_s1_translator:clk, led_s1_translator_avalon_universal_slave_0_agent:clk, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, leftdata:clk, leftdata_s1_translator:clk, leftdata_s1_translator_avalon_universal_slave_0_agent:clk, leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, leftready:clk, leftready_s1_translator:clk, leftready_s1_translator_avalon_universal_slave_0_agent:clk, leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, leftsenddata:clk, leftsenddata_s1_translator:clk, leftsenddata_s1_translator_avalon_universal_slave_0_agent:clk, leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, lrcin:clk, lrcin_s1_translator:clk, lrcin_s1_translator_avalon_universal_slave_0_agent:clk, lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, lrcout:clk, lrcout_s1_translator:clk, lrcout_s1_translator_avalon_universal_slave_0_agent:clk, lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, nios2_qsys:clk, nios2_qsys_data_master_translator:clk, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_instruction_master_translator:clk, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_jtag_debug_module_translator:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2:clk, onchip_memory2_s1_translator:clk, onchip_memory2_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rightdata:clk, rightdata_s1_translator:clk, rightdata_s1_translator_avalon_universal_slave_0_agent:clk, rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rightready:clk, rightready_s1_translator:clk, rightready_s1_translator_avalon_universal_slave_0_agent:clk, rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rightsenddata:clk, rightsenddata_s1_translator:clk, rightsenddata_s1_translator_avalon_universal_slave_0_agent:clk, rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_demux_020:clk, rsp_xbar_demux_021:clk, rsp_xbar_demux_022:clk, rsp_xbar_demux_023:clk, rsp_xbar_demux_024:clk, rsp_xbar_demux_026:clk, rsp_xbar_demux_027:clk, rsp_xbar_demux_028:clk, rsp_xbar_demux_029:clk, rsp_xbar_demux_030:clk, rsp_xbar_demux_031:clk, rsp_xbar_demux_033:clk, rsp_xbar_demux_034:clk, rsp_xbar_demux_035:clk, rsp_xbar_demux_036:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sclk:clk, sclk_s1_translator:clk, sclk_s1_translator_avalon_universal_slave_0_agent:clk, sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sdin:clk, sdin_s1_translator:clk, sdin_s1_translator_avalon_universal_slave_0_agent:clk, sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch0:clk, switch0_s1_translator:clk, switch0_s1_translator_avalon_universal_slave_0_agent:clk, switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch1:clk, switch1_s1_translator:clk, switch1_s1_translator_avalon_universal_slave_0_agent:clk, switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch2:clk, switch2_s1_translator:clk, switch2_s1_translator_avalon_universal_slave_0_agent:clk, switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch3:clk, switch3_s1_translator:clk, switch3_s1_translator_avalon_universal_slave_0_agent:clk, switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch4:clk, switch4_s1_translator:clk, switch4_s1_translator_avalon_universal_slave_0_agent:clk, switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch5:clk, switch5_s1_translator:clk, switch5_s1_translator_avalon_universal_slave_0_agent:clk, switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch6:clk, switch6_s1_translator:clk, switch6_s1_translator_avalon_universal_slave_0_agent:clk, switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch7:clk, switch7_s1_translator:clk, switch7_s1_translator_avalon_universal_slave_0_agent:clk, switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch8:clk, switch8_s1_translator:clk, switch8_s1_translator_avalon_universal_slave_0_agent:clk, switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid_qsys:clock, sysid_qsys_control_slave_translator:clk, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, uart:clk, uart_s1_translator:clk, uart_s1_translator_avalon_universal_slave_0_agent:clk, uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire         nios2_qsys_instruction_master_waitrequest;                                                         // nios2_qsys_instruction_master_translator:av_waitrequest -> nios2_qsys:i_waitrequest
	wire  [19:0] nios2_qsys_instruction_master_address;                                                             // nios2_qsys:i_address -> nios2_qsys_instruction_master_translator:av_address
	wire         nios2_qsys_instruction_master_read;                                                                // nios2_qsys:i_read -> nios2_qsys_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                                                            // nios2_qsys_instruction_master_translator:av_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                                                       // nios2_qsys_instruction_master_translator:av_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         nios2_qsys_data_master_waitrequest;                                                                // nios2_qsys_data_master_translator:av_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                                                                  // nios2_qsys:d_writedata -> nios2_qsys_data_master_translator:av_writedata
	wire  [19:0] nios2_qsys_data_master_address;                                                                    // nios2_qsys:d_address -> nios2_qsys_data_master_translator:av_address
	wire         nios2_qsys_data_master_write;                                                                      // nios2_qsys:d_write -> nios2_qsys_data_master_translator:av_write
	wire         nios2_qsys_data_master_read;                                                                       // nios2_qsys:d_read -> nios2_qsys_data_master_translator:av_read
	wire  [31:0] nios2_qsys_data_master_readdata;                                                                   // nios2_qsys_data_master_translator:av_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                                                                // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_data_master_translator:av_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                                                              // nios2_qsys_data_master_translator:av_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                                                                 // nios2_qsys:d_byteenable -> nios2_qsys_data_master_translator:av_byteenable
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                           // nios2_qsys:jtag_debug_module_waitrequest -> nios2_qsys_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // nios2_qsys_jtag_debug_module_translator:av_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // nios2_qsys_jtag_debug_module_translator:av_address -> nios2_qsys:jtag_debug_module_address
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // nios2_qsys_jtag_debug_module_translator:av_write -> nios2_qsys:jtag_debug_module_write
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read;                                  // nios2_qsys_jtag_debug_module_translator:av_read -> nios2_qsys:jtag_debug_module_read
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // nios2_qsys:jtag_debug_module_readdata -> nios2_qsys_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // nios2_qsys_jtag_debug_module_translator:av_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // nios2_qsys_jtag_debug_module_translator:av_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory2_s1_translator_avalon_anti_slave_0_writedata;                                        // onchip_memory2_s1_translator:av_writedata -> onchip_memory2:writedata
	wire  [15:0] onchip_memory2_s1_translator_avalon_anti_slave_0_address;                                          // onchip_memory2_s1_translator:av_address -> onchip_memory2:address
	wire         onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect;                                       // onchip_memory2_s1_translator:av_chipselect -> onchip_memory2:chipselect
	wire         onchip_memory2_s1_translator_avalon_anti_slave_0_clken;                                            // onchip_memory2_s1_translator:av_clken -> onchip_memory2:clken
	wire         onchip_memory2_s1_translator_avalon_anti_slave_0_write;                                            // onchip_memory2_s1_translator:av_write -> onchip_memory2:write
	wire  [31:0] onchip_memory2_s1_translator_avalon_anti_slave_0_readdata;                                         // onchip_memory2:readdata -> onchip_memory2_s1_translator:av_readdata
	wire   [3:0] onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable;                                       // onchip_memory2_s1_translator:av_byteenable -> onchip_memory2:byteenable
	wire  [15:0] uart_s1_translator_avalon_anti_slave_0_writedata;                                                  // uart_s1_translator:av_writedata -> uart:writedata
	wire   [2:0] uart_s1_translator_avalon_anti_slave_0_address;                                                    // uart_s1_translator:av_address -> uart:address
	wire         uart_s1_translator_avalon_anti_slave_0_chipselect;                                                 // uart_s1_translator:av_chipselect -> uart:chipselect
	wire         uart_s1_translator_avalon_anti_slave_0_write;                                                      // uart_s1_translator:av_write -> uart:write_n
	wire         uart_s1_translator_avalon_anti_slave_0_read;                                                       // uart_s1_translator:av_read -> uart:read_n
	wire  [15:0] uart_s1_translator_avalon_anti_slave_0_readdata;                                                   // uart:readdata -> uart_s1_translator:av_readdata
	wire         uart_s1_translator_avalon_anti_slave_0_begintransfer;                                              // uart_s1_translator:av_begintransfer -> uart:begintransfer
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire   [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [0:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_address;                                   // sysid_qsys_control_slave_translator:av_address -> sysid_qsys:address
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata;                                  // sysid_qsys:readdata -> sysid_qsys_control_slave_translator:av_readdata
	wire  [31:0] led_s1_translator_avalon_anti_slave_0_writedata;                                                   // led_s1_translator:av_writedata -> led:writedata
	wire   [1:0] led_s1_translator_avalon_anti_slave_0_address;                                                     // led_s1_translator:av_address -> led:address
	wire         led_s1_translator_avalon_anti_slave_0_chipselect;                                                  // led_s1_translator:av_chipselect -> led:chipselect
	wire         led_s1_translator_avalon_anti_slave_0_write;                                                       // led_s1_translator:av_write -> led:write_n
	wire  [31:0] led_s1_translator_avalon_anti_slave_0_readdata;                                                    // led:readdata -> led_s1_translator:av_readdata
	wire  [31:0] switch0_s1_translator_avalon_anti_slave_0_writedata;                                               // switch0_s1_translator:av_writedata -> switch0:writedata
	wire   [1:0] switch0_s1_translator_avalon_anti_slave_0_address;                                                 // switch0_s1_translator:av_address -> switch0:address
	wire         switch0_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch0_s1_translator:av_chipselect -> switch0:chipselect
	wire         switch0_s1_translator_avalon_anti_slave_0_write;                                                   // switch0_s1_translator:av_write -> switch0:write_n
	wire  [31:0] switch0_s1_translator_avalon_anti_slave_0_readdata;                                                // switch0:readdata -> switch0_s1_translator:av_readdata
	wire  [31:0] key0_s1_translator_avalon_anti_slave_0_writedata;                                                  // key0_s1_translator:av_writedata -> key0:writedata
	wire   [1:0] key0_s1_translator_avalon_anti_slave_0_address;                                                    // key0_s1_translator:av_address -> key0:address
	wire         key0_s1_translator_avalon_anti_slave_0_chipselect;                                                 // key0_s1_translator:av_chipselect -> key0:chipselect
	wire         key0_s1_translator_avalon_anti_slave_0_write;                                                      // key0_s1_translator:av_write -> key0:write_n
	wire  [31:0] key0_s1_translator_avalon_anti_slave_0_readdata;                                                   // key0:readdata -> key0_s1_translator:av_readdata
	wire   [1:0] adc_s1_translator_avalon_anti_slave_0_address;                                                     // adc_s1_translator:av_address -> adc:address
	wire  [31:0] adc_s1_translator_avalon_anti_slave_0_readdata;                                                    // adc:readdata -> adc_s1_translator:av_readdata
	wire  [31:0] cs_s1_translator_avalon_anti_slave_0_writedata;                                                    // cs_s1_translator:av_writedata -> cs:writedata
	wire   [1:0] cs_s1_translator_avalon_anti_slave_0_address;                                                      // cs_s1_translator:av_address -> cs:address
	wire         cs_s1_translator_avalon_anti_slave_0_chipselect;                                                   // cs_s1_translator:av_chipselect -> cs:chipselect
	wire         cs_s1_translator_avalon_anti_slave_0_write;                                                        // cs_s1_translator:av_write -> cs:write_n
	wire  [31:0] cs_s1_translator_avalon_anti_slave_0_readdata;                                                     // cs:readdata -> cs_s1_translator:av_readdata
	wire  [31:0] sclk_s1_translator_avalon_anti_slave_0_writedata;                                                  // sclk_s1_translator:av_writedata -> sclk:writedata
	wire   [1:0] sclk_s1_translator_avalon_anti_slave_0_address;                                                    // sclk_s1_translator:av_address -> sclk:address
	wire         sclk_s1_translator_avalon_anti_slave_0_chipselect;                                                 // sclk_s1_translator:av_chipselect -> sclk:chipselect
	wire         sclk_s1_translator_avalon_anti_slave_0_write;                                                      // sclk_s1_translator:av_write -> sclk:write_n
	wire  [31:0] sclk_s1_translator_avalon_anti_slave_0_readdata;                                                   // sclk:readdata -> sclk_s1_translator:av_readdata
	wire  [31:0] sdin_s1_translator_avalon_anti_slave_0_writedata;                                                  // sdin_s1_translator:av_writedata -> sdin:writedata
	wire   [1:0] sdin_s1_translator_avalon_anti_slave_0_address;                                                    // sdin_s1_translator:av_address -> sdin:address
	wire         sdin_s1_translator_avalon_anti_slave_0_chipselect;                                                 // sdin_s1_translator:av_chipselect -> sdin:chipselect
	wire         sdin_s1_translator_avalon_anti_slave_0_write;                                                      // sdin_s1_translator:av_write -> sdin:write_n
	wire  [31:0] sdin_s1_translator_avalon_anti_slave_0_readdata;                                                   // sdin:readdata -> sdin_s1_translator:av_readdata
	wire  [31:0] din_s1_translator_avalon_anti_slave_0_writedata;                                                   // din_s1_translator:av_writedata -> din:writedata
	wire   [1:0] din_s1_translator_avalon_anti_slave_0_address;                                                     // din_s1_translator:av_address -> din:address
	wire         din_s1_translator_avalon_anti_slave_0_chipselect;                                                  // din_s1_translator:av_chipselect -> din:chipselect
	wire         din_s1_translator_avalon_anti_slave_0_write;                                                       // din_s1_translator:av_write -> din:write_n
	wire  [31:0] din_s1_translator_avalon_anti_slave_0_readdata;                                                    // din:readdata -> din_s1_translator:av_readdata
	wire  [31:0] bclk_in_s1_translator_avalon_anti_slave_0_writedata;                                               // bclk_in_s1_translator:av_writedata -> bclk_in:writedata
	wire   [1:0] bclk_in_s1_translator_avalon_anti_slave_0_address;                                                 // bclk_in_s1_translator:av_address -> bclk_in:address
	wire         bclk_in_s1_translator_avalon_anti_slave_0_chipselect;                                              // bclk_in_s1_translator:av_chipselect -> bclk_in:chipselect
	wire         bclk_in_s1_translator_avalon_anti_slave_0_write;                                                   // bclk_in_s1_translator:av_write -> bclk_in:write_n
	wire  [31:0] bclk_in_s1_translator_avalon_anti_slave_0_readdata;                                                // bclk_in:readdata -> bclk_in_s1_translator:av_readdata
	wire  [31:0] lrcout_s1_translator_avalon_anti_slave_0_writedata;                                                // lrcout_s1_translator:av_writedata -> lrcout:writedata
	wire   [1:0] lrcout_s1_translator_avalon_anti_slave_0_address;                                                  // lrcout_s1_translator:av_address -> lrcout:address
	wire         lrcout_s1_translator_avalon_anti_slave_0_chipselect;                                               // lrcout_s1_translator:av_chipselect -> lrcout:chipselect
	wire         lrcout_s1_translator_avalon_anti_slave_0_write;                                                    // lrcout_s1_translator:av_write -> lrcout:write_n
	wire  [31:0] lrcout_s1_translator_avalon_anti_slave_0_readdata;                                                 // lrcout:readdata -> lrcout_s1_translator:av_readdata
	wire   [1:0] dout_s1_translator_avalon_anti_slave_0_address;                                                    // dout_s1_translator:av_address -> dout:address
	wire  [31:0] dout_s1_translator_avalon_anti_slave_0_readdata;                                                   // dout:readdata -> dout_s1_translator:av_readdata
	wire  [31:0] bclk_out_s1_translator_avalon_anti_slave_0_writedata;                                              // bclk_out_s1_translator:av_writedata -> bclk_out:writedata
	wire   [1:0] bclk_out_s1_translator_avalon_anti_slave_0_address;                                                // bclk_out_s1_translator:av_address -> bclk_out:address
	wire         bclk_out_s1_translator_avalon_anti_slave_0_chipselect;                                             // bclk_out_s1_translator:av_chipselect -> bclk_out:chipselect
	wire         bclk_out_s1_translator_avalon_anti_slave_0_write;                                                  // bclk_out_s1_translator:av_write -> bclk_out:write_n
	wire  [31:0] bclk_out_s1_translator_avalon_anti_slave_0_readdata;                                               // bclk_out:readdata -> bclk_out_s1_translator:av_readdata
	wire  [31:0] lrcin_s1_translator_avalon_anti_slave_0_writedata;                                                 // lrcin_s1_translator:av_writedata -> lrcin:writedata
	wire   [1:0] lrcin_s1_translator_avalon_anti_slave_0_address;                                                   // lrcin_s1_translator:av_address -> lrcin:address
	wire         lrcin_s1_translator_avalon_anti_slave_0_chipselect;                                                // lrcin_s1_translator:av_chipselect -> lrcin:chipselect
	wire         lrcin_s1_translator_avalon_anti_slave_0_write;                                                     // lrcin_s1_translator:av_write -> lrcin:write_n
	wire  [31:0] lrcin_s1_translator_avalon_anti_slave_0_readdata;                                                  // lrcin:readdata -> lrcin_s1_translator:av_readdata
	wire  [31:0] key1_s1_translator_avalon_anti_slave_0_writedata;                                                  // key1_s1_translator:av_writedata -> key1:writedata
	wire   [1:0] key1_s1_translator_avalon_anti_slave_0_address;                                                    // key1_s1_translator:av_address -> key1:address
	wire         key1_s1_translator_avalon_anti_slave_0_chipselect;                                                 // key1_s1_translator:av_chipselect -> key1:chipselect
	wire         key1_s1_translator_avalon_anti_slave_0_write;                                                      // key1_s1_translator:av_write -> key1:write_n
	wire  [31:0] key1_s1_translator_avalon_anti_slave_0_readdata;                                                   // key1:readdata -> key1_s1_translator:av_readdata
	wire  [31:0] key2_s1_translator_avalon_anti_slave_0_writedata;                                                  // key2_s1_translator:av_writedata -> key2:writedata
	wire   [1:0] key2_s1_translator_avalon_anti_slave_0_address;                                                    // key2_s1_translator:av_address -> key2:address
	wire         key2_s1_translator_avalon_anti_slave_0_chipselect;                                                 // key2_s1_translator:av_chipselect -> key2:chipselect
	wire         key2_s1_translator_avalon_anti_slave_0_write;                                                      // key2_s1_translator:av_write -> key2:write_n
	wire  [31:0] key2_s1_translator_avalon_anti_slave_0_readdata;                                                   // key2:readdata -> key2_s1_translator:av_readdata
	wire  [31:0] key3_s1_translator_avalon_anti_slave_0_writedata;                                                  // key3_s1_translator:av_writedata -> key3:writedata
	wire   [1:0] key3_s1_translator_avalon_anti_slave_0_address;                                                    // key3_s1_translator:av_address -> key3:address
	wire         key3_s1_translator_avalon_anti_slave_0_chipselect;                                                 // key3_s1_translator:av_chipselect -> key3:chipselect
	wire         key3_s1_translator_avalon_anti_slave_0_write;                                                      // key3_s1_translator:av_write -> key3:write_n
	wire  [31:0] key3_s1_translator_avalon_anti_slave_0_readdata;                                                   // key3:readdata -> key3_s1_translator:av_readdata
	wire  [31:0] switch1_s1_translator_avalon_anti_slave_0_writedata;                                               // switch1_s1_translator:av_writedata -> switch1:writedata
	wire   [1:0] switch1_s1_translator_avalon_anti_slave_0_address;                                                 // switch1_s1_translator:av_address -> switch1:address
	wire         switch1_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch1_s1_translator:av_chipselect -> switch1:chipselect
	wire         switch1_s1_translator_avalon_anti_slave_0_write;                                                   // switch1_s1_translator:av_write -> switch1:write_n
	wire  [31:0] switch1_s1_translator_avalon_anti_slave_0_readdata;                                                // switch1:readdata -> switch1_s1_translator:av_readdata
	wire  [31:0] switch2_s1_translator_avalon_anti_slave_0_writedata;                                               // switch2_s1_translator:av_writedata -> switch2:writedata
	wire   [1:0] switch2_s1_translator_avalon_anti_slave_0_address;                                                 // switch2_s1_translator:av_address -> switch2:address
	wire         switch2_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch2_s1_translator:av_chipselect -> switch2:chipselect
	wire         switch2_s1_translator_avalon_anti_slave_0_write;                                                   // switch2_s1_translator:av_write -> switch2:write_n
	wire  [31:0] switch2_s1_translator_avalon_anti_slave_0_readdata;                                                // switch2:readdata -> switch2_s1_translator:av_readdata
	wire  [31:0] switch3_s1_translator_avalon_anti_slave_0_writedata;                                               // switch3_s1_translator:av_writedata -> switch3:writedata
	wire   [1:0] switch3_s1_translator_avalon_anti_slave_0_address;                                                 // switch3_s1_translator:av_address -> switch3:address
	wire         switch3_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch3_s1_translator:av_chipselect -> switch3:chipselect
	wire         switch3_s1_translator_avalon_anti_slave_0_write;                                                   // switch3_s1_translator:av_write -> switch3:write_n
	wire  [31:0] switch3_s1_translator_avalon_anti_slave_0_readdata;                                                // switch3:readdata -> switch3_s1_translator:av_readdata
	wire  [31:0] switch4_s1_translator_avalon_anti_slave_0_writedata;                                               // switch4_s1_translator:av_writedata -> switch4:writedata
	wire   [1:0] switch4_s1_translator_avalon_anti_slave_0_address;                                                 // switch4_s1_translator:av_address -> switch4:address
	wire         switch4_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch4_s1_translator:av_chipselect -> switch4:chipselect
	wire         switch4_s1_translator_avalon_anti_slave_0_write;                                                   // switch4_s1_translator:av_write -> switch4:write_n
	wire  [31:0] switch4_s1_translator_avalon_anti_slave_0_readdata;                                                // switch4:readdata -> switch4_s1_translator:av_readdata
	wire  [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata;                                       // altpll_0_pll_slave_translator:av_writedata -> altpll_0:writedata
	wire   [1:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_address;                                         // altpll_0_pll_slave_translator:av_address -> altpll_0:address
	wire         altpll_0_pll_slave_translator_avalon_anti_slave_0_write;                                           // altpll_0_pll_slave_translator:av_write -> altpll_0:write
	wire         altpll_0_pll_slave_translator_avalon_anti_slave_0_read;                                            // altpll_0_pll_slave_translator:av_read -> altpll_0:read
	wire  [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata;                                        // altpll_0:readdata -> altpll_0_pll_slave_translator:av_readdata
	wire   [1:0] leftdata_s1_translator_avalon_anti_slave_0_address;                                                // leftdata_s1_translator:av_address -> leftdata:address
	wire  [31:0] leftdata_s1_translator_avalon_anti_slave_0_readdata;                                               // leftdata:readdata -> leftdata_s1_translator:av_readdata
	wire   [1:0] rightdata_s1_translator_avalon_anti_slave_0_address;                                               // rightdata_s1_translator:av_address -> rightdata:address
	wire  [31:0] rightdata_s1_translator_avalon_anti_slave_0_readdata;                                              // rightdata:readdata -> rightdata_s1_translator:av_readdata
	wire  [31:0] leftready_s1_translator_avalon_anti_slave_0_writedata;                                             // leftready_s1_translator:av_writedata -> leftready:writedata
	wire   [1:0] leftready_s1_translator_avalon_anti_slave_0_address;                                               // leftready_s1_translator:av_address -> leftready:address
	wire         leftready_s1_translator_avalon_anti_slave_0_chipselect;                                            // leftready_s1_translator:av_chipselect -> leftready:chipselect
	wire         leftready_s1_translator_avalon_anti_slave_0_write;                                                 // leftready_s1_translator:av_write -> leftready:write_n
	wire  [31:0] leftready_s1_translator_avalon_anti_slave_0_readdata;                                              // leftready:readdata -> leftready_s1_translator:av_readdata
	wire  [31:0] rightready_s1_translator_avalon_anti_slave_0_writedata;                                            // rightready_s1_translator:av_writedata -> rightready:writedata
	wire   [1:0] rightready_s1_translator_avalon_anti_slave_0_address;                                              // rightready_s1_translator:av_address -> rightready:address
	wire         rightready_s1_translator_avalon_anti_slave_0_chipselect;                                           // rightready_s1_translator:av_chipselect -> rightready:chipselect
	wire         rightready_s1_translator_avalon_anti_slave_0_write;                                                // rightready_s1_translator:av_write -> rightready:write_n
	wire  [31:0] rightready_s1_translator_avalon_anti_slave_0_readdata;                                             // rightready:readdata -> rightready_s1_translator:av_readdata
	wire  [31:0] leftsenddata_s1_translator_avalon_anti_slave_0_writedata;                                          // leftsenddata_s1_translator:av_writedata -> leftsenddata:writedata
	wire   [1:0] leftsenddata_s1_translator_avalon_anti_slave_0_address;                                            // leftsenddata_s1_translator:av_address -> leftsenddata:address
	wire         leftsenddata_s1_translator_avalon_anti_slave_0_chipselect;                                         // leftsenddata_s1_translator:av_chipselect -> leftsenddata:chipselect
	wire         leftsenddata_s1_translator_avalon_anti_slave_0_write;                                              // leftsenddata_s1_translator:av_write -> leftsenddata:write_n
	wire  [31:0] leftsenddata_s1_translator_avalon_anti_slave_0_readdata;                                           // leftsenddata:readdata -> leftsenddata_s1_translator:av_readdata
	wire  [31:0] rightsenddata_s1_translator_avalon_anti_slave_0_writedata;                                         // rightsenddata_s1_translator:av_writedata -> rightsenddata:writedata
	wire   [1:0] rightsenddata_s1_translator_avalon_anti_slave_0_address;                                           // rightsenddata_s1_translator:av_address -> rightsenddata:address
	wire         rightsenddata_s1_translator_avalon_anti_slave_0_chipselect;                                        // rightsenddata_s1_translator:av_chipselect -> rightsenddata:chipselect
	wire         rightsenddata_s1_translator_avalon_anti_slave_0_write;                                             // rightsenddata_s1_translator:av_write -> rightsenddata:write_n
	wire  [31:0] rightsenddata_s1_translator_avalon_anti_slave_0_readdata;                                          // rightsenddata:readdata -> rightsenddata_s1_translator:av_readdata
	wire  [31:0] clk_12mhz_pll_slave_translator_avalon_anti_slave_0_writedata;                                      // clk_12mhz_pll_slave_translator:av_writedata -> clk_12mhz:writedata
	wire   [1:0] clk_12mhz_pll_slave_translator_avalon_anti_slave_0_address;                                        // clk_12mhz_pll_slave_translator:av_address -> clk_12mhz:address
	wire         clk_12mhz_pll_slave_translator_avalon_anti_slave_0_write;                                          // clk_12mhz_pll_slave_translator:av_write -> clk_12mhz:write
	wire         clk_12mhz_pll_slave_translator_avalon_anti_slave_0_read;                                           // clk_12mhz_pll_slave_translator:av_read -> clk_12mhz:read
	wire  [31:0] clk_12mhz_pll_slave_translator_avalon_anti_slave_0_readdata;                                       // clk_12mhz:readdata -> clk_12mhz_pll_slave_translator:av_readdata
	wire  [31:0] switch5_s1_translator_avalon_anti_slave_0_writedata;                                               // switch5_s1_translator:av_writedata -> switch5:writedata
	wire   [1:0] switch5_s1_translator_avalon_anti_slave_0_address;                                                 // switch5_s1_translator:av_address -> switch5:address
	wire         switch5_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch5_s1_translator:av_chipselect -> switch5:chipselect
	wire         switch5_s1_translator_avalon_anti_slave_0_write;                                                   // switch5_s1_translator:av_write -> switch5:write_n
	wire  [31:0] switch5_s1_translator_avalon_anti_slave_0_readdata;                                                // switch5:readdata -> switch5_s1_translator:av_readdata
	wire  [31:0] switch6_s1_translator_avalon_anti_slave_0_writedata;                                               // switch6_s1_translator:av_writedata -> switch6:writedata
	wire   [1:0] switch6_s1_translator_avalon_anti_slave_0_address;                                                 // switch6_s1_translator:av_address -> switch6:address
	wire         switch6_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch6_s1_translator:av_chipselect -> switch6:chipselect
	wire         switch6_s1_translator_avalon_anti_slave_0_write;                                                   // switch6_s1_translator:av_write -> switch6:write_n
	wire  [31:0] switch6_s1_translator_avalon_anti_slave_0_readdata;                                                // switch6:readdata -> switch6_s1_translator:av_readdata
	wire  [31:0] switch7_s1_translator_avalon_anti_slave_0_writedata;                                               // switch7_s1_translator:av_writedata -> switch7:writedata
	wire   [1:0] switch7_s1_translator_avalon_anti_slave_0_address;                                                 // switch7_s1_translator:av_address -> switch7:address
	wire         switch7_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch7_s1_translator:av_chipselect -> switch7:chipselect
	wire         switch7_s1_translator_avalon_anti_slave_0_write;                                                   // switch7_s1_translator:av_write -> switch7:write_n
	wire  [31:0] switch7_s1_translator_avalon_anti_slave_0_readdata;                                                // switch7:readdata -> switch7_s1_translator:av_readdata
	wire  [31:0] switch8_s1_translator_avalon_anti_slave_0_writedata;                                               // switch8_s1_translator:av_writedata -> switch8:writedata
	wire   [1:0] switch8_s1_translator_avalon_anti_slave_0_address;                                                 // switch8_s1_translator:av_address -> switch8:address
	wire         switch8_s1_translator_avalon_anti_slave_0_chipselect;                                              // switch8_s1_translator:av_chipselect -> switch8:chipselect
	wire         switch8_s1_translator_avalon_anti_slave_0_write;                                                   // switch8_s1_translator:av_write -> switch8:write_n
	wire  [31:0] switch8_s1_translator_avalon_anti_slave_0_readdata;                                                // switch8:readdata -> switch8_s1_translator:av_readdata
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount;                     // nios2_qsys_instruction_master_translator:uav_burstcount -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata;                      // nios2_qsys_instruction_master_translator:uav_writedata -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [19:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_address;                        // nios2_qsys_instruction_master_translator:uav_address -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock;                           // nios2_qsys_instruction_master_translator:uav_lock -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_write;                          // nios2_qsys_instruction_master_translator:uav_write -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_read;                           // nios2_qsys_instruction_master_translator:uav_read -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata;                       // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_instruction_master_translator:uav_readdata
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // nios2_qsys_instruction_master_translator:uav_debugaccess -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable;                     // nios2_qsys_instruction_master_translator:uav_byteenable -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_instruction_master_translator:uav_readdatavalid
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_data_master_translator:uav_burstcount -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_data_master_translator:uav_writedata -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [19:0] nios2_qsys_data_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_data_master_translator:uav_address -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_data_master_translator:uav_lock -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_data_master_translator:uav_write -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_data_master_translator:uav_read -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_data_master_translator:uav_readdata
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_data_master_translator:uav_debugaccess -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_data_master_translator:uav_byteenable -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_data_master_translator:uav_readdatavalid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // nios2_qsys_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_jtag_debug_module_translator:uav_writedata
	wire  [19:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // nios2_qsys_jtag_debug_module_translator:uav_readdata -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // nios2_qsys_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // onchip_memory2_s1_translator:uav_waitrequest -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_s1_translator:uav_writedata
	wire  [19:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_s1_translator:uav_address
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_s1_translator:uav_write
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_s1_translator:uav_lock
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_s1_translator:uav_read
	wire  [31:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // onchip_memory2_s1_translator:uav_readdata -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // onchip_memory2_s1_translator:uav_readdatavalid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_s1_translator:uav_byteenable
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // uart_s1_translator:uav_waitrequest -> uart_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // uart_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_s1_translator:uav_burstcount
	wire  [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // uart_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_s1_translator:uav_writedata
	wire  [19:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // uart_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_s1_translator:uav_address
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // uart_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_s1_translator:uav_write
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // uart_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_s1_translator:uav_lock
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // uart_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_s1_translator:uav_read
	wire  [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // uart_s1_translator:uav_readdata -> uart_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // uart_s1_translator:uav_readdatavalid -> uart_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // uart_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_s1_translator:uav_debugaccess
	wire   [3:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // uart_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_s1_translator:uav_byteenable
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire  [19:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // sysid_qsys_control_slave_translator:uav_waitrequest -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_control_slave_translator:uav_writedata
	wire  [19:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_control_slave_translator:uav_address
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_control_slave_translator:uav_write
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_control_slave_translator:uav_lock
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_control_slave_translator:uav_read
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // sysid_qsys_control_slave_translator:uav_readdata -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // sysid_qsys_control_slave_translator:uav_readdatavalid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_control_slave_translator:uav_byteenable
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // led_s1_translator:uav_waitrequest -> led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_s1_translator:uav_burstcount
	wire  [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_s1_translator:uav_writedata
	wire  [19:0] led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // led_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_s1_translator:uav_address
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // led_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_s1_translator:uav_write
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_s1_translator:uav_lock
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // led_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_s1_translator:uav_read
	wire  [31:0] led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // led_s1_translator:uav_readdata -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // led_s1_translator:uav_readdatavalid -> led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_s1_translator:uav_debugaccess
	wire   [3:0] led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_s1_translator:uav_byteenable
	wire         led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch0_s1_translator:uav_waitrequest -> switch0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch0_s1_translator:uav_burstcount
	wire  [31:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch0_s1_translator:uav_writedata
	wire  [19:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch0_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch0_s1_translator:uav_address
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch0_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch0_s1_translator:uav_write
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch0_s1_translator:uav_lock
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch0_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch0_s1_translator:uav_read
	wire  [31:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch0_s1_translator:uav_readdata -> switch0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch0_s1_translator:uav_readdatavalid -> switch0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch0_s1_translator:uav_debugaccess
	wire   [3:0] switch0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch0_s1_translator:uav_byteenable
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         key0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // key0_s1_translator:uav_waitrequest -> key0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] key0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // key0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key0_s1_translator:uav_burstcount
	wire  [31:0] key0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // key0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key0_s1_translator:uav_writedata
	wire  [19:0] key0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // key0_s1_translator_avalon_universal_slave_0_agent:m0_address -> key0_s1_translator:uav_address
	wire         key0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // key0_s1_translator_avalon_universal_slave_0_agent:m0_write -> key0_s1_translator:uav_write
	wire         key0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // key0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key0_s1_translator:uav_lock
	wire         key0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // key0_s1_translator_avalon_universal_slave_0_agent:m0_read -> key0_s1_translator:uav_read
	wire  [31:0] key0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // key0_s1_translator:uav_readdata -> key0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         key0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // key0_s1_translator:uav_readdatavalid -> key0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         key0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // key0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key0_s1_translator:uav_debugaccess
	wire   [3:0] key0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // key0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key0_s1_translator:uav_byteenable
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // key0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // key0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // key0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] key0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // key0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // key0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // key0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // key0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // key0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         adc_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // adc_s1_translator:uav_waitrequest -> adc_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] adc_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // adc_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> adc_s1_translator:uav_burstcount
	wire  [31:0] adc_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // adc_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> adc_s1_translator:uav_writedata
	wire  [19:0] adc_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // adc_s1_translator_avalon_universal_slave_0_agent:m0_address -> adc_s1_translator:uav_address
	wire         adc_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // adc_s1_translator_avalon_universal_slave_0_agent:m0_write -> adc_s1_translator:uav_write
	wire         adc_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // adc_s1_translator_avalon_universal_slave_0_agent:m0_lock -> adc_s1_translator:uav_lock
	wire         adc_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // adc_s1_translator_avalon_universal_slave_0_agent:m0_read -> adc_s1_translator:uav_read
	wire  [31:0] adc_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // adc_s1_translator:uav_readdata -> adc_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         adc_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // adc_s1_translator:uav_readdatavalid -> adc_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         adc_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // adc_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> adc_s1_translator:uav_debugaccess
	wire   [3:0] adc_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // adc_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> adc_s1_translator:uav_byteenable
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // adc_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // adc_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // adc_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] adc_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // adc_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> adc_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> adc_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> adc_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> adc_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> adc_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // adc_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // adc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> adc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // adc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> adc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // adc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> adc_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // cs_s1_translator:uav_waitrequest -> cs_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] cs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // cs_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> cs_s1_translator:uav_burstcount
	wire  [31:0] cs_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // cs_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> cs_s1_translator:uav_writedata
	wire  [19:0] cs_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // cs_s1_translator_avalon_universal_slave_0_agent:m0_address -> cs_s1_translator:uav_address
	wire         cs_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // cs_s1_translator_avalon_universal_slave_0_agent:m0_write -> cs_s1_translator:uav_write
	wire         cs_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // cs_s1_translator_avalon_universal_slave_0_agent:m0_lock -> cs_s1_translator:uav_lock
	wire         cs_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // cs_s1_translator_avalon_universal_slave_0_agent:m0_read -> cs_s1_translator:uav_read
	wire  [31:0] cs_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // cs_s1_translator:uav_readdata -> cs_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         cs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // cs_s1_translator:uav_readdatavalid -> cs_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         cs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // cs_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cs_s1_translator:uav_debugaccess
	wire   [3:0] cs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // cs_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> cs_s1_translator:uav_byteenable
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // cs_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // cs_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // cs_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] cs_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // cs_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cs_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cs_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cs_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cs_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cs_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // cs_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // cs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // cs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // cs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // sclk_s1_translator:uav_waitrequest -> sclk_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sclk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // sclk_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sclk_s1_translator:uav_burstcount
	wire  [31:0] sclk_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // sclk_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sclk_s1_translator:uav_writedata
	wire  [19:0] sclk_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // sclk_s1_translator_avalon_universal_slave_0_agent:m0_address -> sclk_s1_translator:uav_address
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // sclk_s1_translator_avalon_universal_slave_0_agent:m0_write -> sclk_s1_translator:uav_write
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // sclk_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sclk_s1_translator:uav_lock
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // sclk_s1_translator_avalon_universal_slave_0_agent:m0_read -> sclk_s1_translator:uav_read
	wire  [31:0] sclk_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // sclk_s1_translator:uav_readdata -> sclk_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // sclk_s1_translator:uav_readdatavalid -> sclk_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // sclk_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sclk_s1_translator:uav_debugaccess
	wire   [3:0] sclk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // sclk_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sclk_s1_translator:uav_byteenable
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // sclk_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // sclk_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // sclk_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // sclk_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sclk_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // sclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // sclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // sclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // sclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // sdin_s1_translator:uav_waitrequest -> sdin_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sdin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // sdin_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdin_s1_translator:uav_burstcount
	wire  [31:0] sdin_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // sdin_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdin_s1_translator:uav_writedata
	wire  [19:0] sdin_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // sdin_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdin_s1_translator:uav_address
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // sdin_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdin_s1_translator:uav_write
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // sdin_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdin_s1_translator:uav_lock
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // sdin_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdin_s1_translator:uav_read
	wire  [31:0] sdin_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // sdin_s1_translator:uav_readdata -> sdin_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // sdin_s1_translator:uav_readdatavalid -> sdin_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // sdin_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdin_s1_translator:uav_debugaccess
	wire   [3:0] sdin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // sdin_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdin_s1_translator:uav_byteenable
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // sdin_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // sdin_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // sdin_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // sdin_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdin_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdin_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdin_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdin_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdin_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // sdin_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // sdin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // sdin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // sdin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         din_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // din_s1_translator:uav_waitrequest -> din_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] din_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // din_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> din_s1_translator:uav_burstcount
	wire  [31:0] din_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // din_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> din_s1_translator:uav_writedata
	wire  [19:0] din_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // din_s1_translator_avalon_universal_slave_0_agent:m0_address -> din_s1_translator:uav_address
	wire         din_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // din_s1_translator_avalon_universal_slave_0_agent:m0_write -> din_s1_translator:uav_write
	wire         din_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // din_s1_translator_avalon_universal_slave_0_agent:m0_lock -> din_s1_translator:uav_lock
	wire         din_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // din_s1_translator_avalon_universal_slave_0_agent:m0_read -> din_s1_translator:uav_read
	wire  [31:0] din_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // din_s1_translator:uav_readdata -> din_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         din_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // din_s1_translator:uav_readdatavalid -> din_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         din_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // din_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> din_s1_translator:uav_debugaccess
	wire   [3:0] din_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // din_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> din_s1_translator:uav_byteenable
	wire         din_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // din_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         din_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // din_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         din_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // din_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] din_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // din_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         din_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> din_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> din_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> din_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> din_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> din_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // din_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // din_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> din_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // din_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> din_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // din_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> din_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // bclk_in_s1_translator:uav_waitrequest -> bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> bclk_in_s1_translator:uav_burstcount
	wire  [31:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> bclk_in_s1_translator:uav_writedata
	wire  [19:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_address -> bclk_in_s1_translator:uav_address
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_write -> bclk_in_s1_translator:uav_write
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_lock -> bclk_in_s1_translator:uav_lock
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_read -> bclk_in_s1_translator:uav_read
	wire  [31:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // bclk_in_s1_translator:uav_readdata -> bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // bclk_in_s1_translator:uav_readdatavalid -> bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> bclk_in_s1_translator:uav_debugaccess
	wire   [3:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // bclk_in_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> bclk_in_s1_translator:uav_byteenable
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // bclk_in_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // bclk_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // bclk_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // bclk_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // lrcout_s1_translator:uav_waitrequest -> lrcout_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lrcout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // lrcout_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lrcout_s1_translator:uav_burstcount
	wire  [31:0] lrcout_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // lrcout_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lrcout_s1_translator:uav_writedata
	wire  [19:0] lrcout_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // lrcout_s1_translator_avalon_universal_slave_0_agent:m0_address -> lrcout_s1_translator:uav_address
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // lrcout_s1_translator_avalon_universal_slave_0_agent:m0_write -> lrcout_s1_translator:uav_write
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // lrcout_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lrcout_s1_translator:uav_lock
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // lrcout_s1_translator_avalon_universal_slave_0_agent:m0_read -> lrcout_s1_translator:uav_read
	wire  [31:0] lrcout_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // lrcout_s1_translator:uav_readdata -> lrcout_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // lrcout_s1_translator:uav_readdatavalid -> lrcout_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // lrcout_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lrcout_s1_translator:uav_debugaccess
	wire   [3:0] lrcout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // lrcout_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lrcout_s1_translator:uav_byteenable
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // lrcout_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // lrcout_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // lrcout_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // lrcout_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lrcout_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lrcout_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lrcout_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lrcout_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lrcout_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // lrcout_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // lrcout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lrcout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // lrcout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lrcout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // lrcout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lrcout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         dout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // dout_s1_translator:uav_waitrequest -> dout_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] dout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // dout_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> dout_s1_translator:uav_burstcount
	wire  [31:0] dout_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // dout_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> dout_s1_translator:uav_writedata
	wire  [19:0] dout_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // dout_s1_translator_avalon_universal_slave_0_agent:m0_address -> dout_s1_translator:uav_address
	wire         dout_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // dout_s1_translator_avalon_universal_slave_0_agent:m0_write -> dout_s1_translator:uav_write
	wire         dout_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // dout_s1_translator_avalon_universal_slave_0_agent:m0_lock -> dout_s1_translator:uav_lock
	wire         dout_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // dout_s1_translator_avalon_universal_slave_0_agent:m0_read -> dout_s1_translator:uav_read
	wire  [31:0] dout_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // dout_s1_translator:uav_readdata -> dout_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         dout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // dout_s1_translator:uav_readdatavalid -> dout_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         dout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // dout_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dout_s1_translator:uav_debugaccess
	wire   [3:0] dout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // dout_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> dout_s1_translator:uav_byteenable
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // dout_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // dout_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // dout_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] dout_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // dout_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dout_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dout_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dout_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dout_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dout_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // dout_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // dout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // dout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // dout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dout_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // bclk_out_s1_translator:uav_waitrequest -> bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> bclk_out_s1_translator:uav_burstcount
	wire  [31:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> bclk_out_s1_translator:uav_writedata
	wire  [19:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_address -> bclk_out_s1_translator:uav_address
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_write -> bclk_out_s1_translator:uav_write
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_lock -> bclk_out_s1_translator:uav_lock
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_read -> bclk_out_s1_translator:uav_read
	wire  [31:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // bclk_out_s1_translator:uav_readdata -> bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // bclk_out_s1_translator:uav_readdatavalid -> bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> bclk_out_s1_translator:uav_debugaccess
	wire   [3:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // bclk_out_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> bclk_out_s1_translator:uav_byteenable
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // bclk_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // bclk_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // bclk_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // bclk_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // lrcin_s1_translator:uav_waitrequest -> lrcin_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lrcin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // lrcin_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lrcin_s1_translator:uav_burstcount
	wire  [31:0] lrcin_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // lrcin_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lrcin_s1_translator:uav_writedata
	wire  [19:0] lrcin_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // lrcin_s1_translator_avalon_universal_slave_0_agent:m0_address -> lrcin_s1_translator:uav_address
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // lrcin_s1_translator_avalon_universal_slave_0_agent:m0_write -> lrcin_s1_translator:uav_write
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // lrcin_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lrcin_s1_translator:uav_lock
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // lrcin_s1_translator_avalon_universal_slave_0_agent:m0_read -> lrcin_s1_translator:uav_read
	wire  [31:0] lrcin_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // lrcin_s1_translator:uav_readdata -> lrcin_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // lrcin_s1_translator:uav_readdatavalid -> lrcin_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // lrcin_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lrcin_s1_translator:uav_debugaccess
	wire   [3:0] lrcin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // lrcin_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lrcin_s1_translator:uav_byteenable
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // lrcin_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // lrcin_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // lrcin_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // lrcin_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lrcin_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lrcin_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lrcin_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lrcin_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lrcin_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // lrcin_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // lrcin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lrcin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // lrcin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lrcin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // lrcin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lrcin_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // key1_s1_translator:uav_waitrequest -> key1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // key1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key1_s1_translator:uav_burstcount
	wire  [31:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // key1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key1_s1_translator:uav_writedata
	wire  [19:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // key1_s1_translator_avalon_universal_slave_0_agent:m0_address -> key1_s1_translator:uav_address
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // key1_s1_translator_avalon_universal_slave_0_agent:m0_write -> key1_s1_translator:uav_write
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // key1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key1_s1_translator:uav_lock
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // key1_s1_translator_avalon_universal_slave_0_agent:m0_read -> key1_s1_translator:uav_read
	wire  [31:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // key1_s1_translator:uav_readdata -> key1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // key1_s1_translator:uav_readdatavalid -> key1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         key1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // key1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key1_s1_translator:uav_debugaccess
	wire   [3:0] key1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // key1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key1_s1_translator:uav_byteenable
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // key1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // key1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // key1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] key1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // key1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // key1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // key2_s1_translator:uav_waitrequest -> key2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // key2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key2_s1_translator:uav_burstcount
	wire  [31:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // key2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key2_s1_translator:uav_writedata
	wire  [19:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // key2_s1_translator_avalon_universal_slave_0_agent:m0_address -> key2_s1_translator:uav_address
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // key2_s1_translator_avalon_universal_slave_0_agent:m0_write -> key2_s1_translator:uav_write
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // key2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key2_s1_translator:uav_lock
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // key2_s1_translator_avalon_universal_slave_0_agent:m0_read -> key2_s1_translator:uav_read
	wire  [31:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // key2_s1_translator:uav_readdata -> key2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // key2_s1_translator:uav_readdatavalid -> key2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         key2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // key2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key2_s1_translator:uav_debugaccess
	wire   [3:0] key2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // key2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key2_s1_translator:uav_byteenable
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // key2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // key2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // key2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] key2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // key2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // key2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // key3_s1_translator:uav_waitrequest -> key3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // key3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key3_s1_translator:uav_burstcount
	wire  [31:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // key3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key3_s1_translator:uav_writedata
	wire  [19:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // key3_s1_translator_avalon_universal_slave_0_agent:m0_address -> key3_s1_translator:uav_address
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // key3_s1_translator_avalon_universal_slave_0_agent:m0_write -> key3_s1_translator:uav_write
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // key3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key3_s1_translator:uav_lock
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // key3_s1_translator_avalon_universal_slave_0_agent:m0_read -> key3_s1_translator:uav_read
	wire  [31:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // key3_s1_translator:uav_readdata -> key3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // key3_s1_translator:uav_readdatavalid -> key3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         key3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // key3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key3_s1_translator:uav_debugaccess
	wire   [3:0] key3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // key3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key3_s1_translator:uav_byteenable
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // key3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // key3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // key3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] key3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // key3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // key3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch1_s1_translator:uav_waitrequest -> switch1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch1_s1_translator:uav_burstcount
	wire  [31:0] switch1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch1_s1_translator:uav_writedata
	wire  [19:0] switch1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch1_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch1_s1_translator:uav_address
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch1_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch1_s1_translator:uav_write
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch1_s1_translator:uav_lock
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch1_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch1_s1_translator:uav_read
	wire  [31:0] switch1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch1_s1_translator:uav_readdata -> switch1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch1_s1_translator:uav_readdatavalid -> switch1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch1_s1_translator:uav_debugaccess
	wire   [3:0] switch1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch1_s1_translator:uav_byteenable
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch2_s1_translator:uav_waitrequest -> switch2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch2_s1_translator:uav_burstcount
	wire  [31:0] switch2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch2_s1_translator:uav_writedata
	wire  [19:0] switch2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch2_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch2_s1_translator:uav_address
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch2_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch2_s1_translator:uav_write
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch2_s1_translator:uav_lock
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch2_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch2_s1_translator:uav_read
	wire  [31:0] switch2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch2_s1_translator:uav_readdata -> switch2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch2_s1_translator:uav_readdatavalid -> switch2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch2_s1_translator:uav_debugaccess
	wire   [3:0] switch2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch2_s1_translator:uav_byteenable
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch3_s1_translator:uav_waitrequest -> switch3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch3_s1_translator:uav_burstcount
	wire  [31:0] switch3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch3_s1_translator:uav_writedata
	wire  [19:0] switch3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch3_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch3_s1_translator:uav_address
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch3_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch3_s1_translator:uav_write
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch3_s1_translator:uav_lock
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch3_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch3_s1_translator:uav_read
	wire  [31:0] switch3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch3_s1_translator:uav_readdata -> switch3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch3_s1_translator:uav_readdatavalid -> switch3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch3_s1_translator:uav_debugaccess
	wire   [3:0] switch3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch3_s1_translator:uav_byteenable
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch4_s1_translator:uav_waitrequest -> switch4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch4_s1_translator:uav_burstcount
	wire  [31:0] switch4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch4_s1_translator:uav_writedata
	wire  [19:0] switch4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch4_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch4_s1_translator:uav_address
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch4_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch4_s1_translator:uav_write
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch4_s1_translator:uav_lock
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch4_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch4_s1_translator:uav_read
	wire  [31:0] switch4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch4_s1_translator:uav_readdata -> switch4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch4_s1_translator:uav_readdatavalid -> switch4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch4_s1_translator:uav_debugaccess
	wire   [3:0] switch4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch4_s1_translator:uav_byteenable
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // altpll_0_pll_slave_translator:uav_waitrequest -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> altpll_0_pll_slave_translator:uav_burstcount
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> altpll_0_pll_slave_translator:uav_writedata
	wire  [19:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> altpll_0_pll_slave_translator:uav_address
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> altpll_0_pll_slave_translator:uav_write
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> altpll_0_pll_slave_translator:uav_lock
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> altpll_0_pll_slave_translator:uav_read
	wire  [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // altpll_0_pll_slave_translator:uav_readdata -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // altpll_0_pll_slave_translator:uav_readdatavalid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> altpll_0_pll_slave_translator:uav_debugaccess
	wire   [3:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> altpll_0_pll_slave_translator:uav_byteenable
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [33:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // leftdata_s1_translator:uav_waitrequest -> leftdata_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] leftdata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // leftdata_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> leftdata_s1_translator:uav_burstcount
	wire  [31:0] leftdata_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // leftdata_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> leftdata_s1_translator:uav_writedata
	wire  [19:0] leftdata_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // leftdata_s1_translator_avalon_universal_slave_0_agent:m0_address -> leftdata_s1_translator:uav_address
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // leftdata_s1_translator_avalon_universal_slave_0_agent:m0_write -> leftdata_s1_translator:uav_write
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // leftdata_s1_translator_avalon_universal_slave_0_agent:m0_lock -> leftdata_s1_translator:uav_lock
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // leftdata_s1_translator_avalon_universal_slave_0_agent:m0_read -> leftdata_s1_translator:uav_read
	wire  [31:0] leftdata_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // leftdata_s1_translator:uav_readdata -> leftdata_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // leftdata_s1_translator:uav_readdatavalid -> leftdata_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // leftdata_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> leftdata_s1_translator:uav_debugaccess
	wire   [3:0] leftdata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // leftdata_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> leftdata_s1_translator:uav_byteenable
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // leftdata_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // leftdata_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // leftdata_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // leftdata_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> leftdata_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> leftdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> leftdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> leftdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> leftdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // leftdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // leftdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> leftdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // leftdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> leftdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // leftdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> leftdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // rightdata_s1_translator:uav_waitrequest -> rightdata_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rightdata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // rightdata_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> rightdata_s1_translator:uav_burstcount
	wire  [31:0] rightdata_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // rightdata_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> rightdata_s1_translator:uav_writedata
	wire  [19:0] rightdata_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // rightdata_s1_translator_avalon_universal_slave_0_agent:m0_address -> rightdata_s1_translator:uav_address
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // rightdata_s1_translator_avalon_universal_slave_0_agent:m0_write -> rightdata_s1_translator:uav_write
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // rightdata_s1_translator_avalon_universal_slave_0_agent:m0_lock -> rightdata_s1_translator:uav_lock
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // rightdata_s1_translator_avalon_universal_slave_0_agent:m0_read -> rightdata_s1_translator:uav_read
	wire  [31:0] rightdata_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // rightdata_s1_translator:uav_readdata -> rightdata_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // rightdata_s1_translator:uav_readdatavalid -> rightdata_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // rightdata_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rightdata_s1_translator:uav_debugaccess
	wire   [3:0] rightdata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // rightdata_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> rightdata_s1_translator:uav_byteenable
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // rightdata_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // rightdata_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // rightdata_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // rightdata_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rightdata_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rightdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rightdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rightdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rightdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // rightdata_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // rightdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rightdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // rightdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rightdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // rightdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rightdata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // leftready_s1_translator:uav_waitrequest -> leftready_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] leftready_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // leftready_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> leftready_s1_translator:uav_burstcount
	wire  [31:0] leftready_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // leftready_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> leftready_s1_translator:uav_writedata
	wire  [19:0] leftready_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // leftready_s1_translator_avalon_universal_slave_0_agent:m0_address -> leftready_s1_translator:uav_address
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // leftready_s1_translator_avalon_universal_slave_0_agent:m0_write -> leftready_s1_translator:uav_write
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // leftready_s1_translator_avalon_universal_slave_0_agent:m0_lock -> leftready_s1_translator:uav_lock
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // leftready_s1_translator_avalon_universal_slave_0_agent:m0_read -> leftready_s1_translator:uav_read
	wire  [31:0] leftready_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // leftready_s1_translator:uav_readdata -> leftready_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // leftready_s1_translator:uav_readdatavalid -> leftready_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // leftready_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> leftready_s1_translator:uav_debugaccess
	wire   [3:0] leftready_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // leftready_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> leftready_s1_translator:uav_byteenable
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // leftready_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // leftready_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // leftready_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // leftready_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> leftready_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> leftready_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> leftready_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> leftready_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> leftready_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // leftready_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // leftready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> leftready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // leftready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> leftready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // leftready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> leftready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // rightready_s1_translator:uav_waitrequest -> rightready_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rightready_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // rightready_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> rightready_s1_translator:uav_burstcount
	wire  [31:0] rightready_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // rightready_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> rightready_s1_translator:uav_writedata
	wire  [19:0] rightready_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // rightready_s1_translator_avalon_universal_slave_0_agent:m0_address -> rightready_s1_translator:uav_address
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // rightready_s1_translator_avalon_universal_slave_0_agent:m0_write -> rightready_s1_translator:uav_write
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // rightready_s1_translator_avalon_universal_slave_0_agent:m0_lock -> rightready_s1_translator:uav_lock
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // rightready_s1_translator_avalon_universal_slave_0_agent:m0_read -> rightready_s1_translator:uav_read
	wire  [31:0] rightready_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // rightready_s1_translator:uav_readdata -> rightready_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // rightready_s1_translator:uav_readdatavalid -> rightready_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // rightready_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rightready_s1_translator:uav_debugaccess
	wire   [3:0] rightready_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // rightready_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> rightready_s1_translator:uav_byteenable
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // rightready_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // rightready_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // rightready_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // rightready_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rightready_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rightready_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rightready_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rightready_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rightready_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // rightready_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // rightready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rightready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // rightready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rightready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // rightready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rightready_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // leftsenddata_s1_translator:uav_waitrequest -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> leftsenddata_s1_translator:uav_burstcount
	wire  [31:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> leftsenddata_s1_translator:uav_writedata
	wire  [19:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_address -> leftsenddata_s1_translator:uav_address
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_write -> leftsenddata_s1_translator:uav_write
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_lock -> leftsenddata_s1_translator:uav_lock
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_read -> leftsenddata_s1_translator:uav_read
	wire  [31:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // leftsenddata_s1_translator:uav_readdata -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // leftsenddata_s1_translator:uav_readdatavalid -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> leftsenddata_s1_translator:uav_debugaccess
	wire   [3:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // leftsenddata_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> leftsenddata_s1_translator:uav_byteenable
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // rightsenddata_s1_translator:uav_waitrequest -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> rightsenddata_s1_translator:uav_burstcount
	wire  [31:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                           // rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> rightsenddata_s1_translator:uav_writedata
	wire  [19:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_address;                             // rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_address -> rightsenddata_s1_translator:uav_address
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_write;                               // rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_write -> rightsenddata_s1_translator:uav_write
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                // rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_lock -> rightsenddata_s1_translator:uav_lock
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_read;                                // rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_read -> rightsenddata_s1_translator:uav_read
	wire  [31:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                            // rightsenddata_s1_translator:uav_readdata -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // rightsenddata_s1_translator:uav_readdatavalid -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rightsenddata_s1_translator:uav_debugaccess
	wire   [3:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // rightsenddata_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> rightsenddata_s1_translator:uav_byteenable
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                         // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // clk_12mhz_pll_slave_translator:uav_waitrequest -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> clk_12mhz_pll_slave_translator:uav_burstcount
	wire  [31:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> clk_12mhz_pll_slave_translator:uav_writedata
	wire  [19:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> clk_12mhz_pll_slave_translator:uav_address
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> clk_12mhz_pll_slave_translator:uav_write
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> clk_12mhz_pll_slave_translator:uav_lock
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> clk_12mhz_pll_slave_translator:uav_read
	wire  [31:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // clk_12mhz_pll_slave_translator:uav_readdata -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // clk_12mhz_pll_slave_translator:uav_readdatavalid -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> clk_12mhz_pll_slave_translator:uav_debugaccess
	wire   [3:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> clk_12mhz_pll_slave_translator:uav_byteenable
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [33:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch5_s1_translator:uav_waitrequest -> switch5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch5_s1_translator:uav_burstcount
	wire  [31:0] switch5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch5_s1_translator:uav_writedata
	wire  [19:0] switch5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch5_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch5_s1_translator:uav_address
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch5_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch5_s1_translator:uav_write
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch5_s1_translator:uav_lock
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch5_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch5_s1_translator:uav_read
	wire  [31:0] switch5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch5_s1_translator:uav_readdata -> switch5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch5_s1_translator:uav_readdatavalid -> switch5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch5_s1_translator:uav_debugaccess
	wire   [3:0] switch5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch5_s1_translator:uav_byteenable
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch6_s1_translator:uav_waitrequest -> switch6_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch6_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch6_s1_translator:uav_burstcount
	wire  [31:0] switch6_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch6_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch6_s1_translator:uav_writedata
	wire  [19:0] switch6_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch6_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch6_s1_translator:uav_address
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch6_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch6_s1_translator:uav_write
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch6_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch6_s1_translator:uav_lock
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch6_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch6_s1_translator:uav_read
	wire  [31:0] switch6_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch6_s1_translator:uav_readdata -> switch6_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch6_s1_translator:uav_readdatavalid -> switch6_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch6_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch6_s1_translator:uav_debugaccess
	wire   [3:0] switch6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch6_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch6_s1_translator:uav_byteenable
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch6_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch6_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch6_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch6_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch6_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch6_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch6_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch6_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch6_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch6_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch7_s1_translator:uav_waitrequest -> switch7_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch7_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch7_s1_translator:uav_burstcount
	wire  [31:0] switch7_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch7_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch7_s1_translator:uav_writedata
	wire  [19:0] switch7_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch7_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch7_s1_translator:uav_address
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch7_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch7_s1_translator:uav_write
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch7_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch7_s1_translator:uav_lock
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch7_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch7_s1_translator:uav_read
	wire  [31:0] switch7_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch7_s1_translator:uav_readdata -> switch7_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch7_s1_translator:uav_readdatavalid -> switch7_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch7_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch7_s1_translator:uav_debugaccess
	wire   [3:0] switch7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch7_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch7_s1_translator:uav_byteenable
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch7_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch7_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch7_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch7_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch7_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch7_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch7_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch7_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch7_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch7_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // switch8_s1_translator:uav_waitrequest -> switch8_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch8_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // switch8_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch8_s1_translator:uav_burstcount
	wire  [31:0] switch8_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // switch8_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch8_s1_translator:uav_writedata
	wire  [19:0] switch8_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // switch8_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch8_s1_translator:uav_address
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // switch8_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch8_s1_translator:uav_write
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // switch8_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch8_s1_translator:uav_lock
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // switch8_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch8_s1_translator:uav_read
	wire  [31:0] switch8_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // switch8_s1_translator:uav_readdata -> switch8_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // switch8_s1_translator:uav_readdatavalid -> switch8_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // switch8_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch8_s1_translator:uav_debugaccess
	wire   [3:0] switch8_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // switch8_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch8_s1_translator:uav_byteenable
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // switch8_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // switch8_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // switch8_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [99:0] switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // switch8_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch8_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch8_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch8_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch8_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [99:0] switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch8_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // switch8_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // switch8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // switch8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // switch8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch8_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [98:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [98:0] nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [98:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [98:0] onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_001:sink_ready -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // uart_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // uart_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // uart_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [98:0] uart_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // uart_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_002:sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [98:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_003:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [98:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_004:sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [98:0] led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_005:sink_ready -> led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [98:0] switch0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         switch0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_006:sink_ready -> switch0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // key0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // key0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // key0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [98:0] key0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // key0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         key0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_007:sink_ready -> key0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // adc_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // adc_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // adc_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [98:0] adc_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // adc_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         adc_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_008:sink_ready -> adc_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // cs_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // cs_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // cs_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [98:0] cs_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // cs_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         cs_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_009:sink_ready -> cs_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // sclk_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // sclk_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // sclk_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [98:0] sclk_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // sclk_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         sclk_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_010:sink_ready -> sclk_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // sdin_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // sdin_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // sdin_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [98:0] sdin_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // sdin_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         sdin_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_011:sink_ready -> sdin_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         din_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // din_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         din_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // din_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         din_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // din_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [98:0] din_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // din_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         din_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_012:sink_ready -> din_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // bclk_in_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // bclk_in_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // bclk_in_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [98:0] bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // bclk_in_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_013:sink_ready -> bclk_in_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // lrcout_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // lrcout_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // lrcout_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [98:0] lrcout_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // lrcout_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         lrcout_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_014:sink_ready -> lrcout_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // dout_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // dout_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // dout_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [98:0] dout_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // dout_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         dout_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_015:sink_ready -> dout_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // bclk_out_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // bclk_out_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // bclk_out_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [98:0] bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // bclk_out_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_016:sink_ready -> bclk_out_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // lrcin_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // lrcin_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // lrcin_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [98:0] lrcin_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // lrcin_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire         lrcin_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_017:sink_ready -> lrcin_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // key1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // key1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // key1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [98:0] key1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // key1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire         key1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_018:sink_ready -> key1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // key2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // key2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // key2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [98:0] key2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // key2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire         key2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_019:sink_ready -> key2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // key3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // key3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // key3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [98:0] key3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // key3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire         key3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_020:sink_ready -> key3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [98:0] switch1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire         switch1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_021:sink_ready -> switch1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [98:0] switch2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire         switch2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_022:sink_ready -> switch2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [98:0] switch3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire         switch3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_023:sink_ready -> switch3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [98:0] switch4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire         switch4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_024:sink_ready -> switch4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [98:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire         altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_025:sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // leftdata_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // leftdata_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // leftdata_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire  [98:0] leftdata_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // leftdata_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire         leftdata_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_026:sink_ready -> leftdata_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // rightdata_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // rightdata_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // rightdata_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire  [98:0] rightdata_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // rightdata_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire         rightdata_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_027:sink_ready -> rightdata_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // leftready_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // leftready_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // leftready_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire  [98:0] leftready_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // leftready_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire         leftready_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_028:sink_ready -> leftready_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // rightready_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // rightready_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // rightready_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire  [98:0] rightready_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // rightready_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire         rightready_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_029:sink_ready -> rightready_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire  [98:0] leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // leftsenddata_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire         leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_030:sink_ready -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_valid;                               // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire  [98:0] rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_data;                                // rightsenddata_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire         rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_031:sink_ready -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire  [98:0] clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire         clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_032:sink_ready -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_033:sink_endofpacket
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_033:sink_valid
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_033:sink_startofpacket
	wire  [98:0] switch5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_033:sink_data
	wire         switch5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_033:sink_ready -> switch5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch6_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_034:sink_endofpacket
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch6_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_034:sink_valid
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch6_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_034:sink_startofpacket
	wire  [98:0] switch6_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch6_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_034:sink_data
	wire         switch6_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_034:sink_ready -> switch6_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch7_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_035:sink_endofpacket
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch7_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_035:sink_valid
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch7_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_035:sink_startofpacket
	wire  [98:0] switch7_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch7_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_035:sink_data
	wire         switch7_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_035:sink_ready -> switch7_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // switch8_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_036:sink_endofpacket
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // switch8_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_036:sink_valid
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // switch8_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_036:sink_startofpacket
	wire  [98:0] switch8_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // switch8_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_036:sink_data
	wire         switch8_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_036:sink_ready -> switch8_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                       // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                             // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                     // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [98:0] addr_router_src_data;                                                                              // addr_router:src_data -> limiter:cmd_sink_data
	wire  [36:0] addr_router_src_channel;                                                                           // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                             // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                       // limiter:rsp_src_endofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                             // limiter:rsp_src_valid -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                     // limiter:rsp_src_startofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [98:0] limiter_rsp_src_data;                                                                              // limiter:rsp_src_data -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [36:0] limiter_rsp_src_channel;                                                                           // limiter:rsp_src_channel -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                             // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                   // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                         // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                 // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [98:0] addr_router_001_src_data;                                                                          // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire  [36:0] addr_router_001_src_channel;                                                                       // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                         // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                   // limiter_001:rsp_src_endofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                         // limiter_001:rsp_src_valid -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                 // limiter_001:rsp_src_startofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [98:0] limiter_001_rsp_src_data;                                                                          // limiter_001:rsp_src_data -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [36:0] limiter_001_rsp_src_channel;                                                                       // limiter_001:rsp_src_channel -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         rst_controller_reset_out_reset;                                                                    // rst_controller:reset_out -> [adc:reset_n, adc_s1_translator:reset, adc_s1_translator_avalon_universal_slave_0_agent:reset, adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, bclk_in:reset_n, bclk_in_s1_translator:reset, bclk_in_s1_translator_avalon_universal_slave_0_agent:reset, bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, bclk_out:reset_n, bclk_out_s1_translator:reset, bclk_out_s1_translator_avalon_universal_slave_0_agent:reset, bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:out_reset, crosser_003:out_reset, cs:reset_n, cs_s1_translator:reset, cs_s1_translator_avalon_universal_slave_0_agent:reset, cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, din:reset_n, din_s1_translator:reset, din_s1_translator_avalon_universal_slave_0_agent:reset, din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dout:reset_n, dout_s1_translator:reset, dout_s1_translator_avalon_universal_slave_0_agent:reset, dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, id_router_030:reset, id_router_031:reset, id_router_033:reset, id_router_034:reset, id_router_035:reset, id_router_036:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key0:reset_n, key0_s1_translator:reset, key0_s1_translator_avalon_universal_slave_0_agent:reset, key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key1:reset_n, key1_s1_translator:reset, key1_s1_translator_avalon_universal_slave_0_agent:reset, key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key2:reset_n, key2_s1_translator:reset, key2_s1_translator_avalon_universal_slave_0_agent:reset, key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key3:reset_n, key3_s1_translator:reset, key3_s1_translator_avalon_universal_slave_0_agent:reset, key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led:reset_n, led_s1_translator:reset, led_s1_translator_avalon_universal_slave_0_agent:reset, led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, leftdata:reset_n, leftdata_s1_translator:reset, leftdata_s1_translator_avalon_universal_slave_0_agent:reset, leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, leftready:reset_n, leftready_s1_translator:reset, leftready_s1_translator_avalon_universal_slave_0_agent:reset, leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, leftsenddata:reset_n, leftsenddata_s1_translator:reset, leftsenddata_s1_translator_avalon_universal_slave_0_agent:reset, leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, lrcin:reset_n, lrcin_s1_translator:reset, lrcin_s1_translator_avalon_universal_slave_0_agent:reset, lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lrcout:reset_n, lrcout_s1_translator:reset, lrcout_s1_translator_avalon_universal_slave_0_agent:reset, lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys:reset_n, nios2_qsys_data_master_translator:reset, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_instruction_master_translator:reset, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_jtag_debug_module_translator:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2:reset, onchip_memory2_s1_translator:reset, onchip_memory2_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rightdata:reset_n, rightdata_s1_translator:reset, rightdata_s1_translator_avalon_universal_slave_0_agent:reset, rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rightready:reset_n, rightready_s1_translator:reset, rightready_s1_translator_avalon_universal_slave_0_agent:reset, rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rightsenddata:reset_n, rightsenddata_s1_translator:reset, rightsenddata_s1_translator_avalon_universal_slave_0_agent:reset, rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_031:reset, rsp_xbar_demux_033:reset, rsp_xbar_demux_034:reset, rsp_xbar_demux_035:reset, rsp_xbar_demux_036:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sclk:reset_n, sclk_s1_translator:reset, sclk_s1_translator_avalon_universal_slave_0_agent:reset, sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sdin:reset_n, sdin_s1_translator:reset, sdin_s1_translator_avalon_universal_slave_0_agent:reset, sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch0:reset_n, switch0_s1_translator:reset, switch0_s1_translator_avalon_universal_slave_0_agent:reset, switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch1:reset_n, switch1_s1_translator:reset, switch1_s1_translator_avalon_universal_slave_0_agent:reset, switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch2:reset_n, switch2_s1_translator:reset, switch2_s1_translator_avalon_universal_slave_0_agent:reset, switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch3:reset_n, switch3_s1_translator:reset, switch3_s1_translator_avalon_universal_slave_0_agent:reset, switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch4:reset_n, switch4_s1_translator:reset, switch4_s1_translator_avalon_universal_slave_0_agent:reset, switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch5:reset_n, switch5_s1_translator:reset, switch5_s1_translator_avalon_universal_slave_0_agent:reset, switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch6:reset_n, switch6_s1_translator:reset, switch6_s1_translator_avalon_universal_slave_0_agent:reset, switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch7:reset_n, switch7_s1_translator:reset, switch7_s1_translator_avalon_universal_slave_0_agent:reset, switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch8:reset_n, switch8_s1_translator:reset, switch8_s1_translator_avalon_universal_slave_0_agent:reset, switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys:reset_n, sysid_qsys_control_slave_translator:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart:reset_n, uart_s1_translator:reset, uart_s1_translator_avalon_universal_slave_0_agent:reset, uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_reset_out_reset_req;                                                                // rst_controller:reset_req -> onchip_memory2:reset_req
	wire         nios2_qsys_jtag_debug_module_reset_reset;                                                          // nios2_qsys:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                                                // rst_controller_001:reset_out -> [altpll_0:reset, altpll_0_pll_slave_translator:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, clk_12mhz:reset, clk_12mhz_pll_slave_translator:reset, clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:reset, clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:in_reset, id_router_025:reset, id_router_032:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_032:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                   // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                         // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                 // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src0_data;                                                                          // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [36:0] cmd_xbar_demux_src0_channel;                                                                       // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                         // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                   // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                         // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                 // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [98:0] cmd_xbar_demux_src1_data;                                                                          // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [36:0] cmd_xbar_demux_src1_channel;                                                                       // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                         // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                               // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                     // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                             // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src0_data;                                                                      // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [36:0] cmd_xbar_demux_001_src0_channel;                                                                   // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                     // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                               // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                     // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                             // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src1_data;                                                                      // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [36:0] cmd_xbar_demux_001_src1_channel;                                                                   // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                     // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                               // cmd_xbar_demux_001:src2_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                     // cmd_xbar_demux_001:src2_valid -> uart_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                             // cmd_xbar_demux_001:src2_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src2_data;                                                                      // cmd_xbar_demux_001:src2_data -> uart_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src2_channel;                                                                   // cmd_xbar_demux_001:src2_channel -> uart_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                               // cmd_xbar_demux_001:src3_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                     // cmd_xbar_demux_001:src3_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                             // cmd_xbar_demux_001:src3_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src3_data;                                                                      // cmd_xbar_demux_001:src3_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src3_channel;                                                                   // cmd_xbar_demux_001:src3_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                               // cmd_xbar_demux_001:src4_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                     // cmd_xbar_demux_001:src4_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                             // cmd_xbar_demux_001:src4_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src4_data;                                                                      // cmd_xbar_demux_001:src4_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src4_channel;                                                                   // cmd_xbar_demux_001:src4_channel -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                               // cmd_xbar_demux_001:src5_endofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                     // cmd_xbar_demux_001:src5_valid -> led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                             // cmd_xbar_demux_001:src5_startofpacket -> led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src5_data;                                                                      // cmd_xbar_demux_001:src5_data -> led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src5_channel;                                                                   // cmd_xbar_demux_001:src5_channel -> led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                               // cmd_xbar_demux_001:src6_endofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                     // cmd_xbar_demux_001:src6_valid -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                             // cmd_xbar_demux_001:src6_startofpacket -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src6_data;                                                                      // cmd_xbar_demux_001:src6_data -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src6_channel;                                                                   // cmd_xbar_demux_001:src6_channel -> switch0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                               // cmd_xbar_demux_001:src7_endofpacket -> key0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                     // cmd_xbar_demux_001:src7_valid -> key0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                             // cmd_xbar_demux_001:src7_startofpacket -> key0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src7_data;                                                                      // cmd_xbar_demux_001:src7_data -> key0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src7_channel;                                                                   // cmd_xbar_demux_001:src7_channel -> key0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                               // cmd_xbar_demux_001:src8_endofpacket -> adc_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                     // cmd_xbar_demux_001:src8_valid -> adc_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                             // cmd_xbar_demux_001:src8_startofpacket -> adc_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src8_data;                                                                      // cmd_xbar_demux_001:src8_data -> adc_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src8_channel;                                                                   // cmd_xbar_demux_001:src8_channel -> adc_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                               // cmd_xbar_demux_001:src9_endofpacket -> cs_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                     // cmd_xbar_demux_001:src9_valid -> cs_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                             // cmd_xbar_demux_001:src9_startofpacket -> cs_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src9_data;                                                                      // cmd_xbar_demux_001:src9_data -> cs_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src9_channel;                                                                   // cmd_xbar_demux_001:src9_channel -> cs_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                              // cmd_xbar_demux_001:src10_endofpacket -> sclk_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                    // cmd_xbar_demux_001:src10_valid -> sclk_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                            // cmd_xbar_demux_001:src10_startofpacket -> sclk_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src10_data;                                                                     // cmd_xbar_demux_001:src10_data -> sclk_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src10_channel;                                                                  // cmd_xbar_demux_001:src10_channel -> sclk_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                              // cmd_xbar_demux_001:src11_endofpacket -> sdin_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                    // cmd_xbar_demux_001:src11_valid -> sdin_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                            // cmd_xbar_demux_001:src11_startofpacket -> sdin_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src11_data;                                                                     // cmd_xbar_demux_001:src11_data -> sdin_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src11_channel;                                                                  // cmd_xbar_demux_001:src11_channel -> sdin_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                              // cmd_xbar_demux_001:src12_endofpacket -> din_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                    // cmd_xbar_demux_001:src12_valid -> din_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                            // cmd_xbar_demux_001:src12_startofpacket -> din_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src12_data;                                                                     // cmd_xbar_demux_001:src12_data -> din_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src12_channel;                                                                  // cmd_xbar_demux_001:src12_channel -> din_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src13_endofpacket;                                                              // cmd_xbar_demux_001:src13_endofpacket -> bclk_in_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src13_valid;                                                                    // cmd_xbar_demux_001:src13_valid -> bclk_in_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src13_startofpacket;                                                            // cmd_xbar_demux_001:src13_startofpacket -> bclk_in_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src13_data;                                                                     // cmd_xbar_demux_001:src13_data -> bclk_in_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src13_channel;                                                                  // cmd_xbar_demux_001:src13_channel -> bclk_in_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src14_endofpacket;                                                              // cmd_xbar_demux_001:src14_endofpacket -> lrcout_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src14_valid;                                                                    // cmd_xbar_demux_001:src14_valid -> lrcout_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src14_startofpacket;                                                            // cmd_xbar_demux_001:src14_startofpacket -> lrcout_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src14_data;                                                                     // cmd_xbar_demux_001:src14_data -> lrcout_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src14_channel;                                                                  // cmd_xbar_demux_001:src14_channel -> lrcout_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src15_endofpacket;                                                              // cmd_xbar_demux_001:src15_endofpacket -> dout_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src15_valid;                                                                    // cmd_xbar_demux_001:src15_valid -> dout_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src15_startofpacket;                                                            // cmd_xbar_demux_001:src15_startofpacket -> dout_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src15_data;                                                                     // cmd_xbar_demux_001:src15_data -> dout_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src15_channel;                                                                  // cmd_xbar_demux_001:src15_channel -> dout_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src16_endofpacket;                                                              // cmd_xbar_demux_001:src16_endofpacket -> bclk_out_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src16_valid;                                                                    // cmd_xbar_demux_001:src16_valid -> bclk_out_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src16_startofpacket;                                                            // cmd_xbar_demux_001:src16_startofpacket -> bclk_out_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src16_data;                                                                     // cmd_xbar_demux_001:src16_data -> bclk_out_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src16_channel;                                                                  // cmd_xbar_demux_001:src16_channel -> bclk_out_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src17_endofpacket;                                                              // cmd_xbar_demux_001:src17_endofpacket -> lrcin_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src17_valid;                                                                    // cmd_xbar_demux_001:src17_valid -> lrcin_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src17_startofpacket;                                                            // cmd_xbar_demux_001:src17_startofpacket -> lrcin_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src17_data;                                                                     // cmd_xbar_demux_001:src17_data -> lrcin_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src17_channel;                                                                  // cmd_xbar_demux_001:src17_channel -> lrcin_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src18_endofpacket;                                                              // cmd_xbar_demux_001:src18_endofpacket -> key1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src18_valid;                                                                    // cmd_xbar_demux_001:src18_valid -> key1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src18_startofpacket;                                                            // cmd_xbar_demux_001:src18_startofpacket -> key1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src18_data;                                                                     // cmd_xbar_demux_001:src18_data -> key1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src18_channel;                                                                  // cmd_xbar_demux_001:src18_channel -> key1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src19_endofpacket;                                                              // cmd_xbar_demux_001:src19_endofpacket -> key2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src19_valid;                                                                    // cmd_xbar_demux_001:src19_valid -> key2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src19_startofpacket;                                                            // cmd_xbar_demux_001:src19_startofpacket -> key2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src19_data;                                                                     // cmd_xbar_demux_001:src19_data -> key2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src19_channel;                                                                  // cmd_xbar_demux_001:src19_channel -> key2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src20_endofpacket;                                                              // cmd_xbar_demux_001:src20_endofpacket -> key3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src20_valid;                                                                    // cmd_xbar_demux_001:src20_valid -> key3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src20_startofpacket;                                                            // cmd_xbar_demux_001:src20_startofpacket -> key3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src20_data;                                                                     // cmd_xbar_demux_001:src20_data -> key3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src20_channel;                                                                  // cmd_xbar_demux_001:src20_channel -> key3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src21_endofpacket;                                                              // cmd_xbar_demux_001:src21_endofpacket -> switch1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src21_valid;                                                                    // cmd_xbar_demux_001:src21_valid -> switch1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src21_startofpacket;                                                            // cmd_xbar_demux_001:src21_startofpacket -> switch1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src21_data;                                                                     // cmd_xbar_demux_001:src21_data -> switch1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src21_channel;                                                                  // cmd_xbar_demux_001:src21_channel -> switch1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src22_endofpacket;                                                              // cmd_xbar_demux_001:src22_endofpacket -> switch2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src22_valid;                                                                    // cmd_xbar_demux_001:src22_valid -> switch2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src22_startofpacket;                                                            // cmd_xbar_demux_001:src22_startofpacket -> switch2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src22_data;                                                                     // cmd_xbar_demux_001:src22_data -> switch2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src22_channel;                                                                  // cmd_xbar_demux_001:src22_channel -> switch2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src23_endofpacket;                                                              // cmd_xbar_demux_001:src23_endofpacket -> switch3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src23_valid;                                                                    // cmd_xbar_demux_001:src23_valid -> switch3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src23_startofpacket;                                                            // cmd_xbar_demux_001:src23_startofpacket -> switch3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src23_data;                                                                     // cmd_xbar_demux_001:src23_data -> switch3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src23_channel;                                                                  // cmd_xbar_demux_001:src23_channel -> switch3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src24_endofpacket;                                                              // cmd_xbar_demux_001:src24_endofpacket -> switch4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src24_valid;                                                                    // cmd_xbar_demux_001:src24_valid -> switch4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src24_startofpacket;                                                            // cmd_xbar_demux_001:src24_startofpacket -> switch4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src24_data;                                                                     // cmd_xbar_demux_001:src24_data -> switch4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src24_channel;                                                                  // cmd_xbar_demux_001:src24_channel -> switch4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src26_endofpacket;                                                              // cmd_xbar_demux_001:src26_endofpacket -> leftdata_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src26_valid;                                                                    // cmd_xbar_demux_001:src26_valid -> leftdata_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src26_startofpacket;                                                            // cmd_xbar_demux_001:src26_startofpacket -> leftdata_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src26_data;                                                                     // cmd_xbar_demux_001:src26_data -> leftdata_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src26_channel;                                                                  // cmd_xbar_demux_001:src26_channel -> leftdata_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src27_endofpacket;                                                              // cmd_xbar_demux_001:src27_endofpacket -> rightdata_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src27_valid;                                                                    // cmd_xbar_demux_001:src27_valid -> rightdata_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src27_startofpacket;                                                            // cmd_xbar_demux_001:src27_startofpacket -> rightdata_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src27_data;                                                                     // cmd_xbar_demux_001:src27_data -> rightdata_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src27_channel;                                                                  // cmd_xbar_demux_001:src27_channel -> rightdata_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src28_endofpacket;                                                              // cmd_xbar_demux_001:src28_endofpacket -> leftready_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src28_valid;                                                                    // cmd_xbar_demux_001:src28_valid -> leftready_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src28_startofpacket;                                                            // cmd_xbar_demux_001:src28_startofpacket -> leftready_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src28_data;                                                                     // cmd_xbar_demux_001:src28_data -> leftready_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src28_channel;                                                                  // cmd_xbar_demux_001:src28_channel -> leftready_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src29_endofpacket;                                                              // cmd_xbar_demux_001:src29_endofpacket -> rightready_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src29_valid;                                                                    // cmd_xbar_demux_001:src29_valid -> rightready_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src29_startofpacket;                                                            // cmd_xbar_demux_001:src29_startofpacket -> rightready_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src29_data;                                                                     // cmd_xbar_demux_001:src29_data -> rightready_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src29_channel;                                                                  // cmd_xbar_demux_001:src29_channel -> rightready_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src30_endofpacket;                                                              // cmd_xbar_demux_001:src30_endofpacket -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src30_valid;                                                                    // cmd_xbar_demux_001:src30_valid -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src30_startofpacket;                                                            // cmd_xbar_demux_001:src30_startofpacket -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src30_data;                                                                     // cmd_xbar_demux_001:src30_data -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src30_channel;                                                                  // cmd_xbar_demux_001:src30_channel -> leftsenddata_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src31_endofpacket;                                                              // cmd_xbar_demux_001:src31_endofpacket -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src31_valid;                                                                    // cmd_xbar_demux_001:src31_valid -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src31_startofpacket;                                                            // cmd_xbar_demux_001:src31_startofpacket -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src31_data;                                                                     // cmd_xbar_demux_001:src31_data -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src31_channel;                                                                  // cmd_xbar_demux_001:src31_channel -> rightsenddata_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src33_endofpacket;                                                              // cmd_xbar_demux_001:src33_endofpacket -> switch5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src33_valid;                                                                    // cmd_xbar_demux_001:src33_valid -> switch5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src33_startofpacket;                                                            // cmd_xbar_demux_001:src33_startofpacket -> switch5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src33_data;                                                                     // cmd_xbar_demux_001:src33_data -> switch5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src33_channel;                                                                  // cmd_xbar_demux_001:src33_channel -> switch5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src34_endofpacket;                                                              // cmd_xbar_demux_001:src34_endofpacket -> switch6_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src34_valid;                                                                    // cmd_xbar_demux_001:src34_valid -> switch6_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src34_startofpacket;                                                            // cmd_xbar_demux_001:src34_startofpacket -> switch6_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src34_data;                                                                     // cmd_xbar_demux_001:src34_data -> switch6_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src34_channel;                                                                  // cmd_xbar_demux_001:src34_channel -> switch6_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src35_endofpacket;                                                              // cmd_xbar_demux_001:src35_endofpacket -> switch7_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src35_valid;                                                                    // cmd_xbar_demux_001:src35_valid -> switch7_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src35_startofpacket;                                                            // cmd_xbar_demux_001:src35_startofpacket -> switch7_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src35_data;                                                                     // cmd_xbar_demux_001:src35_data -> switch7_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src35_channel;                                                                  // cmd_xbar_demux_001:src35_channel -> switch7_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src36_endofpacket;                                                              // cmd_xbar_demux_001:src36_endofpacket -> switch8_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src36_valid;                                                                    // cmd_xbar_demux_001:src36_valid -> switch8_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src36_startofpacket;                                                            // cmd_xbar_demux_001:src36_startofpacket -> switch8_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src36_data;                                                                     // cmd_xbar_demux_001:src36_data -> switch8_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_demux_001_src36_channel;                                                                  // cmd_xbar_demux_001:src36_channel -> switch8_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                   // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                         // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                 // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [98:0] rsp_xbar_demux_src0_data;                                                                          // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [36:0] rsp_xbar_demux_src0_channel;                                                                       // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                         // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                   // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                         // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                 // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [98:0] rsp_xbar_demux_src1_data;                                                                          // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [36:0] rsp_xbar_demux_src1_channel;                                                                       // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                         // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                               // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                     // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                             // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [98:0] rsp_xbar_demux_001_src0_data;                                                                      // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [36:0] rsp_xbar_demux_001_src0_channel;                                                                   // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                     // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                               // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                     // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                             // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [98:0] rsp_xbar_demux_001_src1_data;                                                                      // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [36:0] rsp_xbar_demux_001_src1_channel;                                                                   // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                     // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                               // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                     // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                             // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [98:0] rsp_xbar_demux_002_src0_data;                                                                      // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire  [36:0] rsp_xbar_demux_002_src0_channel;                                                                   // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                     // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                               // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                     // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                             // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [98:0] rsp_xbar_demux_003_src0_data;                                                                      // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire  [36:0] rsp_xbar_demux_003_src0_channel;                                                                   // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                     // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                               // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                     // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                             // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [98:0] rsp_xbar_demux_004_src0_data;                                                                      // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire  [36:0] rsp_xbar_demux_004_src0_channel;                                                                   // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                     // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                               // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                     // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                             // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [98:0] rsp_xbar_demux_005_src0_data;                                                                      // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [36:0] rsp_xbar_demux_005_src0_channel;                                                                   // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                     // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                               // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                     // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                             // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [98:0] rsp_xbar_demux_006_src0_data;                                                                      // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [36:0] rsp_xbar_demux_006_src0_channel;                                                                   // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                     // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                               // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                     // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                             // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [98:0] rsp_xbar_demux_007_src0_data;                                                                      // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [36:0] rsp_xbar_demux_007_src0_channel;                                                                   // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                     // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                               // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                     // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                             // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [98:0] rsp_xbar_demux_008_src0_data;                                                                      // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [36:0] rsp_xbar_demux_008_src0_channel;                                                                   // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                     // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                               // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                     // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                             // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [98:0] rsp_xbar_demux_009_src0_data;                                                                      // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [36:0] rsp_xbar_demux_009_src0_channel;                                                                   // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                     // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                               // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                     // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                             // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [98:0] rsp_xbar_demux_010_src0_data;                                                                      // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [36:0] rsp_xbar_demux_010_src0_channel;                                                                   // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                     // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                               // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                     // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                             // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [98:0] rsp_xbar_demux_011_src0_data;                                                                      // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire  [36:0] rsp_xbar_demux_011_src0_channel;                                                                   // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                     // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                               // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                     // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                             // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [98:0] rsp_xbar_demux_012_src0_data;                                                                      // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire  [36:0] rsp_xbar_demux_012_src0_channel;                                                                   // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                     // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                               // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                     // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                             // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [98:0] rsp_xbar_demux_013_src0_data;                                                                      // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire  [36:0] rsp_xbar_demux_013_src0_channel;                                                                   // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                     // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                               // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                                     // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                             // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [98:0] rsp_xbar_demux_014_src0_data;                                                                      // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire  [36:0] rsp_xbar_demux_014_src0_channel;                                                                   // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                                     // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                               // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                                     // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                             // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [98:0] rsp_xbar_demux_015_src0_data;                                                                      // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire  [36:0] rsp_xbar_demux_015_src0_channel;                                                                   // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                                     // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                               // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                                     // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                             // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [98:0] rsp_xbar_demux_016_src0_data;                                                                      // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire  [36:0] rsp_xbar_demux_016_src0_channel;                                                                   // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                                     // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire         rsp_xbar_demux_017_src0_endofpacket;                                                               // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire         rsp_xbar_demux_017_src0_valid;                                                                     // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire         rsp_xbar_demux_017_src0_startofpacket;                                                             // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [98:0] rsp_xbar_demux_017_src0_data;                                                                      // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire  [36:0] rsp_xbar_demux_017_src0_channel;                                                                   // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire         rsp_xbar_demux_017_src0_ready;                                                                     // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire         rsp_xbar_demux_018_src0_endofpacket;                                                               // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire         rsp_xbar_demux_018_src0_valid;                                                                     // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire         rsp_xbar_demux_018_src0_startofpacket;                                                             // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [98:0] rsp_xbar_demux_018_src0_data;                                                                      // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire  [36:0] rsp_xbar_demux_018_src0_channel;                                                                   // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire         rsp_xbar_demux_018_src0_ready;                                                                     // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire         rsp_xbar_demux_019_src0_endofpacket;                                                               // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire         rsp_xbar_demux_019_src0_valid;                                                                     // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire         rsp_xbar_demux_019_src0_startofpacket;                                                             // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [98:0] rsp_xbar_demux_019_src0_data;                                                                      // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire  [36:0] rsp_xbar_demux_019_src0_channel;                                                                   // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire         rsp_xbar_demux_019_src0_ready;                                                                     // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire         rsp_xbar_demux_020_src0_endofpacket;                                                               // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire         rsp_xbar_demux_020_src0_valid;                                                                     // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	wire         rsp_xbar_demux_020_src0_startofpacket;                                                             // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [98:0] rsp_xbar_demux_020_src0_data;                                                                      // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	wire  [36:0] rsp_xbar_demux_020_src0_channel;                                                                   // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	wire         rsp_xbar_demux_020_src0_ready;                                                                     // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire         rsp_xbar_demux_021_src0_endofpacket;                                                               // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire         rsp_xbar_demux_021_src0_valid;                                                                     // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	wire         rsp_xbar_demux_021_src0_startofpacket;                                                             // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [98:0] rsp_xbar_demux_021_src0_data;                                                                      // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	wire  [36:0] rsp_xbar_demux_021_src0_channel;                                                                   // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	wire         rsp_xbar_demux_021_src0_ready;                                                                     // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire         rsp_xbar_demux_022_src0_endofpacket;                                                               // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire         rsp_xbar_demux_022_src0_valid;                                                                     // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	wire         rsp_xbar_demux_022_src0_startofpacket;                                                             // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [98:0] rsp_xbar_demux_022_src0_data;                                                                      // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	wire  [36:0] rsp_xbar_demux_022_src0_channel;                                                                   // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	wire         rsp_xbar_demux_022_src0_ready;                                                                     // rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire         rsp_xbar_demux_023_src0_endofpacket;                                                               // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink23_endofpacket
	wire         rsp_xbar_demux_023_src0_valid;                                                                     // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink23_valid
	wire         rsp_xbar_demux_023_src0_startofpacket;                                                             // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink23_startofpacket
	wire  [98:0] rsp_xbar_demux_023_src0_data;                                                                      // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink23_data
	wire  [36:0] rsp_xbar_demux_023_src0_channel;                                                                   // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink23_channel
	wire         rsp_xbar_demux_023_src0_ready;                                                                     // rsp_xbar_mux_001:sink23_ready -> rsp_xbar_demux_023:src0_ready
	wire         rsp_xbar_demux_024_src0_endofpacket;                                                               // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink24_endofpacket
	wire         rsp_xbar_demux_024_src0_valid;                                                                     // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink24_valid
	wire         rsp_xbar_demux_024_src0_startofpacket;                                                             // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink24_startofpacket
	wire  [98:0] rsp_xbar_demux_024_src0_data;                                                                      // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink24_data
	wire  [36:0] rsp_xbar_demux_024_src0_channel;                                                                   // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink24_channel
	wire         rsp_xbar_demux_024_src0_ready;                                                                     // rsp_xbar_mux_001:sink24_ready -> rsp_xbar_demux_024:src0_ready
	wire         rsp_xbar_demux_026_src0_endofpacket;                                                               // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_001:sink26_endofpacket
	wire         rsp_xbar_demux_026_src0_valid;                                                                     // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_001:sink26_valid
	wire         rsp_xbar_demux_026_src0_startofpacket;                                                             // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_001:sink26_startofpacket
	wire  [98:0] rsp_xbar_demux_026_src0_data;                                                                      // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_001:sink26_data
	wire  [36:0] rsp_xbar_demux_026_src0_channel;                                                                   // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_001:sink26_channel
	wire         rsp_xbar_demux_026_src0_ready;                                                                     // rsp_xbar_mux_001:sink26_ready -> rsp_xbar_demux_026:src0_ready
	wire         rsp_xbar_demux_027_src0_endofpacket;                                                               // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_001:sink27_endofpacket
	wire         rsp_xbar_demux_027_src0_valid;                                                                     // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_001:sink27_valid
	wire         rsp_xbar_demux_027_src0_startofpacket;                                                             // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_001:sink27_startofpacket
	wire  [98:0] rsp_xbar_demux_027_src0_data;                                                                      // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_001:sink27_data
	wire  [36:0] rsp_xbar_demux_027_src0_channel;                                                                   // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_001:sink27_channel
	wire         rsp_xbar_demux_027_src0_ready;                                                                     // rsp_xbar_mux_001:sink27_ready -> rsp_xbar_demux_027:src0_ready
	wire         rsp_xbar_demux_028_src0_endofpacket;                                                               // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_001:sink28_endofpacket
	wire         rsp_xbar_demux_028_src0_valid;                                                                     // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_001:sink28_valid
	wire         rsp_xbar_demux_028_src0_startofpacket;                                                             // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_001:sink28_startofpacket
	wire  [98:0] rsp_xbar_demux_028_src0_data;                                                                      // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_001:sink28_data
	wire  [36:0] rsp_xbar_demux_028_src0_channel;                                                                   // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_001:sink28_channel
	wire         rsp_xbar_demux_028_src0_ready;                                                                     // rsp_xbar_mux_001:sink28_ready -> rsp_xbar_demux_028:src0_ready
	wire         rsp_xbar_demux_029_src0_endofpacket;                                                               // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_001:sink29_endofpacket
	wire         rsp_xbar_demux_029_src0_valid;                                                                     // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_001:sink29_valid
	wire         rsp_xbar_demux_029_src0_startofpacket;                                                             // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_001:sink29_startofpacket
	wire  [98:0] rsp_xbar_demux_029_src0_data;                                                                      // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_001:sink29_data
	wire  [36:0] rsp_xbar_demux_029_src0_channel;                                                                   // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_001:sink29_channel
	wire         rsp_xbar_demux_029_src0_ready;                                                                     // rsp_xbar_mux_001:sink29_ready -> rsp_xbar_demux_029:src0_ready
	wire         rsp_xbar_demux_030_src0_endofpacket;                                                               // rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux_001:sink30_endofpacket
	wire         rsp_xbar_demux_030_src0_valid;                                                                     // rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux_001:sink30_valid
	wire         rsp_xbar_demux_030_src0_startofpacket;                                                             // rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux_001:sink30_startofpacket
	wire  [98:0] rsp_xbar_demux_030_src0_data;                                                                      // rsp_xbar_demux_030:src0_data -> rsp_xbar_mux_001:sink30_data
	wire  [36:0] rsp_xbar_demux_030_src0_channel;                                                                   // rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux_001:sink30_channel
	wire         rsp_xbar_demux_030_src0_ready;                                                                     // rsp_xbar_mux_001:sink30_ready -> rsp_xbar_demux_030:src0_ready
	wire         rsp_xbar_demux_031_src0_endofpacket;                                                               // rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux_001:sink31_endofpacket
	wire         rsp_xbar_demux_031_src0_valid;                                                                     // rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux_001:sink31_valid
	wire         rsp_xbar_demux_031_src0_startofpacket;                                                             // rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux_001:sink31_startofpacket
	wire  [98:0] rsp_xbar_demux_031_src0_data;                                                                      // rsp_xbar_demux_031:src0_data -> rsp_xbar_mux_001:sink31_data
	wire  [36:0] rsp_xbar_demux_031_src0_channel;                                                                   // rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux_001:sink31_channel
	wire         rsp_xbar_demux_031_src0_ready;                                                                     // rsp_xbar_mux_001:sink31_ready -> rsp_xbar_demux_031:src0_ready
	wire         rsp_xbar_demux_033_src0_endofpacket;                                                               // rsp_xbar_demux_033:src0_endofpacket -> rsp_xbar_mux_001:sink33_endofpacket
	wire         rsp_xbar_demux_033_src0_valid;                                                                     // rsp_xbar_demux_033:src0_valid -> rsp_xbar_mux_001:sink33_valid
	wire         rsp_xbar_demux_033_src0_startofpacket;                                                             // rsp_xbar_demux_033:src0_startofpacket -> rsp_xbar_mux_001:sink33_startofpacket
	wire  [98:0] rsp_xbar_demux_033_src0_data;                                                                      // rsp_xbar_demux_033:src0_data -> rsp_xbar_mux_001:sink33_data
	wire  [36:0] rsp_xbar_demux_033_src0_channel;                                                                   // rsp_xbar_demux_033:src0_channel -> rsp_xbar_mux_001:sink33_channel
	wire         rsp_xbar_demux_033_src0_ready;                                                                     // rsp_xbar_mux_001:sink33_ready -> rsp_xbar_demux_033:src0_ready
	wire         rsp_xbar_demux_034_src0_endofpacket;                                                               // rsp_xbar_demux_034:src0_endofpacket -> rsp_xbar_mux_001:sink34_endofpacket
	wire         rsp_xbar_demux_034_src0_valid;                                                                     // rsp_xbar_demux_034:src0_valid -> rsp_xbar_mux_001:sink34_valid
	wire         rsp_xbar_demux_034_src0_startofpacket;                                                             // rsp_xbar_demux_034:src0_startofpacket -> rsp_xbar_mux_001:sink34_startofpacket
	wire  [98:0] rsp_xbar_demux_034_src0_data;                                                                      // rsp_xbar_demux_034:src0_data -> rsp_xbar_mux_001:sink34_data
	wire  [36:0] rsp_xbar_demux_034_src0_channel;                                                                   // rsp_xbar_demux_034:src0_channel -> rsp_xbar_mux_001:sink34_channel
	wire         rsp_xbar_demux_034_src0_ready;                                                                     // rsp_xbar_mux_001:sink34_ready -> rsp_xbar_demux_034:src0_ready
	wire         rsp_xbar_demux_035_src0_endofpacket;                                                               // rsp_xbar_demux_035:src0_endofpacket -> rsp_xbar_mux_001:sink35_endofpacket
	wire         rsp_xbar_demux_035_src0_valid;                                                                     // rsp_xbar_demux_035:src0_valid -> rsp_xbar_mux_001:sink35_valid
	wire         rsp_xbar_demux_035_src0_startofpacket;                                                             // rsp_xbar_demux_035:src0_startofpacket -> rsp_xbar_mux_001:sink35_startofpacket
	wire  [98:0] rsp_xbar_demux_035_src0_data;                                                                      // rsp_xbar_demux_035:src0_data -> rsp_xbar_mux_001:sink35_data
	wire  [36:0] rsp_xbar_demux_035_src0_channel;                                                                   // rsp_xbar_demux_035:src0_channel -> rsp_xbar_mux_001:sink35_channel
	wire         rsp_xbar_demux_035_src0_ready;                                                                     // rsp_xbar_mux_001:sink35_ready -> rsp_xbar_demux_035:src0_ready
	wire         rsp_xbar_demux_036_src0_endofpacket;                                                               // rsp_xbar_demux_036:src0_endofpacket -> rsp_xbar_mux_001:sink36_endofpacket
	wire         rsp_xbar_demux_036_src0_valid;                                                                     // rsp_xbar_demux_036:src0_valid -> rsp_xbar_mux_001:sink36_valid
	wire         rsp_xbar_demux_036_src0_startofpacket;                                                             // rsp_xbar_demux_036:src0_startofpacket -> rsp_xbar_mux_001:sink36_startofpacket
	wire  [98:0] rsp_xbar_demux_036_src0_data;                                                                      // rsp_xbar_demux_036:src0_data -> rsp_xbar_mux_001:sink36_data
	wire  [36:0] rsp_xbar_demux_036_src0_channel;                                                                   // rsp_xbar_demux_036:src0_channel -> rsp_xbar_mux_001:sink36_channel
	wire         rsp_xbar_demux_036_src0_ready;                                                                     // rsp_xbar_mux_001:sink36_ready -> rsp_xbar_demux_036:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                       // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                     // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [98:0] limiter_cmd_src_data;                                                                              // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [36:0] limiter_cmd_src_channel;                                                                           // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                             // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                      // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                            // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                    // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [98:0] rsp_xbar_mux_src_data;                                                                             // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [36:0] rsp_xbar_mux_src_channel;                                                                          // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                            // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                   // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                 // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [98:0] limiter_001_cmd_src_data;                                                                          // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire  [36:0] limiter_001_cmd_src_channel;                                                                       // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                         // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                  // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                        // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [98:0] rsp_xbar_mux_001_src_data;                                                                         // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire  [36:0] rsp_xbar_mux_001_src_channel;                                                                      // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                        // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                      // cmd_xbar_mux:src_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                            // cmd_xbar_mux:src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                    // cmd_xbar_mux:src_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_src_data;                                                                             // cmd_xbar_mux:src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_mux_src_channel;                                                                          // cmd_xbar_mux:src_channel -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                         // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                               // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                       // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [98:0] id_router_src_data;                                                                                // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [36:0] id_router_src_channel;                                                                             // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                               // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                  // cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                        // cmd_xbar_mux_001:src_valid -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                // cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] cmd_xbar_mux_001_src_data;                                                                         // cmd_xbar_mux_001:src_data -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] cmd_xbar_mux_001_src_channel;                                                                      // cmd_xbar_mux_001:src_channel -> onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                        // onchip_memory2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                     // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                           // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                   // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [98:0] id_router_001_src_data;                                                                            // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [36:0] id_router_001_src_channel;                                                                         // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                           // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_001_src2_ready;                                                                     // uart_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire         id_router_002_src_endofpacket;                                                                     // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                           // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                   // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [98:0] id_router_002_src_data;                                                                            // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [36:0] id_router_002_src_channel;                                                                         // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                           // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                     // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                           // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                   // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [98:0] id_router_003_src_data;                                                                            // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [36:0] id_router_003_src_channel;                                                                         // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                           // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                     // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                           // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                   // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [98:0] id_router_004_src_data;                                                                            // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [36:0] id_router_004_src_channel;                                                                         // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                           // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                     // led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                     // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                           // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                   // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [98:0] id_router_005_src_data;                                                                            // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [36:0] id_router_005_src_channel;                                                                         // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                           // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                     // switch0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                     // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                           // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                   // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [98:0] id_router_006_src_data;                                                                            // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [36:0] id_router_006_src_channel;                                                                         // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                           // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                     // key0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                     // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                           // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                   // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [98:0] id_router_007_src_data;                                                                            // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [36:0] id_router_007_src_channel;                                                                         // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                           // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                     // adc_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                     // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                           // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                   // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [98:0] id_router_008_src_data;                                                                            // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [36:0] id_router_008_src_channel;                                                                         // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                           // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_demux_001_src9_ready;                                                                     // cs_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire         id_router_009_src_endofpacket;                                                                     // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                           // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                   // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [98:0] id_router_009_src_data;                                                                            // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [36:0] id_router_009_src_channel;                                                                         // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                           // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_demux_001_src10_ready;                                                                    // sclk_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire         id_router_010_src_endofpacket;                                                                     // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                           // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                   // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [98:0] id_router_010_src_data;                                                                            // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [36:0] id_router_010_src_channel;                                                                         // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                           // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_001_src11_ready;                                                                    // sdin_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire         id_router_011_src_endofpacket;                                                                     // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                           // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                   // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [98:0] id_router_011_src_data;                                                                            // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [36:0] id_router_011_src_channel;                                                                         // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                           // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_demux_001_src12_ready;                                                                    // din_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire         id_router_012_src_endofpacket;                                                                     // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                           // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                   // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [98:0] id_router_012_src_data;                                                                            // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [36:0] id_router_012_src_channel;                                                                         // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                           // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_demux_001_src13_ready;                                                                    // bclk_in_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire         id_router_013_src_endofpacket;                                                                     // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                           // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                   // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [98:0] id_router_013_src_data;                                                                            // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [36:0] id_router_013_src_channel;                                                                         // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                           // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_demux_001_src14_ready;                                                                    // lrcout_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire         id_router_014_src_endofpacket;                                                                     // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         id_router_014_src_valid;                                                                           // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire         id_router_014_src_startofpacket;                                                                   // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [98:0] id_router_014_src_data;                                                                            // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire  [36:0] id_router_014_src_channel;                                                                         // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire         id_router_014_src_ready;                                                                           // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire         cmd_xbar_demux_001_src15_ready;                                                                    // dout_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire         id_router_015_src_endofpacket;                                                                     // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         id_router_015_src_valid;                                                                           // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire         id_router_015_src_startofpacket;                                                                   // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [98:0] id_router_015_src_data;                                                                            // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire  [36:0] id_router_015_src_channel;                                                                         // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire         id_router_015_src_ready;                                                                           // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire         cmd_xbar_demux_001_src16_ready;                                                                    // bclk_out_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire         id_router_016_src_endofpacket;                                                                     // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         id_router_016_src_valid;                                                                           // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire         id_router_016_src_startofpacket;                                                                   // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [98:0] id_router_016_src_data;                                                                            // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire  [36:0] id_router_016_src_channel;                                                                         // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire         id_router_016_src_ready;                                                                           // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire         cmd_xbar_demux_001_src17_ready;                                                                    // lrcin_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire         id_router_017_src_endofpacket;                                                                     // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire         id_router_017_src_valid;                                                                           // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire         id_router_017_src_startofpacket;                                                                   // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [98:0] id_router_017_src_data;                                                                            // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire  [36:0] id_router_017_src_channel;                                                                         // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire         id_router_017_src_ready;                                                                           // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire         cmd_xbar_demux_001_src18_ready;                                                                    // key1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire         id_router_018_src_endofpacket;                                                                     // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire         id_router_018_src_valid;                                                                           // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire         id_router_018_src_startofpacket;                                                                   // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [98:0] id_router_018_src_data;                                                                            // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire  [36:0] id_router_018_src_channel;                                                                         // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire         id_router_018_src_ready;                                                                           // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire         cmd_xbar_demux_001_src19_ready;                                                                    // key2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	wire         id_router_019_src_endofpacket;                                                                     // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire         id_router_019_src_valid;                                                                           // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire         id_router_019_src_startofpacket;                                                                   // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [98:0] id_router_019_src_data;                                                                            // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire  [36:0] id_router_019_src_channel;                                                                         // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire         id_router_019_src_ready;                                                                           // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire         cmd_xbar_demux_001_src20_ready;                                                                    // key3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	wire         id_router_020_src_endofpacket;                                                                     // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire         id_router_020_src_valid;                                                                           // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire         id_router_020_src_startofpacket;                                                                   // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [98:0] id_router_020_src_data;                                                                            // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire  [36:0] id_router_020_src_channel;                                                                         // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire         id_router_020_src_ready;                                                                           // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire         cmd_xbar_demux_001_src21_ready;                                                                    // switch1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src21_ready
	wire         id_router_021_src_endofpacket;                                                                     // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire         id_router_021_src_valid;                                                                           // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire         id_router_021_src_startofpacket;                                                                   // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [98:0] id_router_021_src_data;                                                                            // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire  [36:0] id_router_021_src_channel;                                                                         // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire         id_router_021_src_ready;                                                                           // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire         cmd_xbar_demux_001_src22_ready;                                                                    // switch2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	wire         id_router_022_src_endofpacket;                                                                     // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire         id_router_022_src_valid;                                                                           // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire         id_router_022_src_startofpacket;                                                                   // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [98:0] id_router_022_src_data;                                                                            // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire  [36:0] id_router_022_src_channel;                                                                         // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire         id_router_022_src_ready;                                                                           // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire         cmd_xbar_demux_001_src23_ready;                                                                    // switch3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src23_ready
	wire         id_router_023_src_endofpacket;                                                                     // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire         id_router_023_src_valid;                                                                           // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire         id_router_023_src_startofpacket;                                                                   // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [98:0] id_router_023_src_data;                                                                            // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire  [36:0] id_router_023_src_channel;                                                                         // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire         id_router_023_src_ready;                                                                           // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire         cmd_xbar_demux_001_src24_ready;                                                                    // switch4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src24_ready
	wire         id_router_024_src_endofpacket;                                                                     // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire         id_router_024_src_valid;                                                                           // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire         id_router_024_src_startofpacket;                                                                   // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [98:0] id_router_024_src_data;                                                                            // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire  [36:0] id_router_024_src_channel;                                                                         // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire         id_router_024_src_ready;                                                                           // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire         crosser_out_ready;                                                                                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire         id_router_025_src_endofpacket;                                                                     // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire         id_router_025_src_valid;                                                                           // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire         id_router_025_src_startofpacket;                                                                   // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [98:0] id_router_025_src_data;                                                                            // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire  [36:0] id_router_025_src_channel;                                                                         // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire         id_router_025_src_ready;                                                                           // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire         cmd_xbar_demux_001_src26_ready;                                                                    // leftdata_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src26_ready
	wire         id_router_026_src_endofpacket;                                                                     // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire         id_router_026_src_valid;                                                                           // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire         id_router_026_src_startofpacket;                                                                   // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire  [98:0] id_router_026_src_data;                                                                            // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire  [36:0] id_router_026_src_channel;                                                                         // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire         id_router_026_src_ready;                                                                           // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire         cmd_xbar_demux_001_src27_ready;                                                                    // rightdata_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src27_ready
	wire         id_router_027_src_endofpacket;                                                                     // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire         id_router_027_src_valid;                                                                           // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire         id_router_027_src_startofpacket;                                                                   // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire  [98:0] id_router_027_src_data;                                                                            // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire  [36:0] id_router_027_src_channel;                                                                         // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire         id_router_027_src_ready;                                                                           // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire         cmd_xbar_demux_001_src28_ready;                                                                    // leftready_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src28_ready
	wire         id_router_028_src_endofpacket;                                                                     // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire         id_router_028_src_valid;                                                                           // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire         id_router_028_src_startofpacket;                                                                   // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire  [98:0] id_router_028_src_data;                                                                            // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire  [36:0] id_router_028_src_channel;                                                                         // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire         id_router_028_src_ready;                                                                           // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire         cmd_xbar_demux_001_src29_ready;                                                                    // rightready_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src29_ready
	wire         id_router_029_src_endofpacket;                                                                     // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire         id_router_029_src_valid;                                                                           // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire         id_router_029_src_startofpacket;                                                                   // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire  [98:0] id_router_029_src_data;                                                                            // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire  [36:0] id_router_029_src_channel;                                                                         // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire         id_router_029_src_ready;                                                                           // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire         cmd_xbar_demux_001_src30_ready;                                                                    // leftsenddata_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src30_ready
	wire         id_router_030_src_endofpacket;                                                                     // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire         id_router_030_src_valid;                                                                           // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire         id_router_030_src_startofpacket;                                                                   // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire  [98:0] id_router_030_src_data;                                                                            // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire  [36:0] id_router_030_src_channel;                                                                         // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire         id_router_030_src_ready;                                                                           // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire         cmd_xbar_demux_001_src31_ready;                                                                    // rightsenddata_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src31_ready
	wire         id_router_031_src_endofpacket;                                                                     // id_router_031:src_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire         id_router_031_src_valid;                                                                           // id_router_031:src_valid -> rsp_xbar_demux_031:sink_valid
	wire         id_router_031_src_startofpacket;                                                                   // id_router_031:src_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire  [98:0] id_router_031_src_data;                                                                            // id_router_031:src_data -> rsp_xbar_demux_031:sink_data
	wire  [36:0] id_router_031_src_channel;                                                                         // id_router_031:src_channel -> rsp_xbar_demux_031:sink_channel
	wire         id_router_031_src_ready;                                                                           // rsp_xbar_demux_031:sink_ready -> id_router_031:src_ready
	wire         crosser_001_out_ready;                                                                             // clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	wire         id_router_032_src_endofpacket;                                                                     // id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire         id_router_032_src_valid;                                                                           // id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	wire         id_router_032_src_startofpacket;                                                                   // id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire  [98:0] id_router_032_src_data;                                                                            // id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	wire  [36:0] id_router_032_src_channel;                                                                         // id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	wire         id_router_032_src_ready;                                                                           // rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	wire         cmd_xbar_demux_001_src33_ready;                                                                    // switch5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src33_ready
	wire         id_router_033_src_endofpacket;                                                                     // id_router_033:src_endofpacket -> rsp_xbar_demux_033:sink_endofpacket
	wire         id_router_033_src_valid;                                                                           // id_router_033:src_valid -> rsp_xbar_demux_033:sink_valid
	wire         id_router_033_src_startofpacket;                                                                   // id_router_033:src_startofpacket -> rsp_xbar_demux_033:sink_startofpacket
	wire  [98:0] id_router_033_src_data;                                                                            // id_router_033:src_data -> rsp_xbar_demux_033:sink_data
	wire  [36:0] id_router_033_src_channel;                                                                         // id_router_033:src_channel -> rsp_xbar_demux_033:sink_channel
	wire         id_router_033_src_ready;                                                                           // rsp_xbar_demux_033:sink_ready -> id_router_033:src_ready
	wire         cmd_xbar_demux_001_src34_ready;                                                                    // switch6_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src34_ready
	wire         id_router_034_src_endofpacket;                                                                     // id_router_034:src_endofpacket -> rsp_xbar_demux_034:sink_endofpacket
	wire         id_router_034_src_valid;                                                                           // id_router_034:src_valid -> rsp_xbar_demux_034:sink_valid
	wire         id_router_034_src_startofpacket;                                                                   // id_router_034:src_startofpacket -> rsp_xbar_demux_034:sink_startofpacket
	wire  [98:0] id_router_034_src_data;                                                                            // id_router_034:src_data -> rsp_xbar_demux_034:sink_data
	wire  [36:0] id_router_034_src_channel;                                                                         // id_router_034:src_channel -> rsp_xbar_demux_034:sink_channel
	wire         id_router_034_src_ready;                                                                           // rsp_xbar_demux_034:sink_ready -> id_router_034:src_ready
	wire         cmd_xbar_demux_001_src35_ready;                                                                    // switch7_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src35_ready
	wire         id_router_035_src_endofpacket;                                                                     // id_router_035:src_endofpacket -> rsp_xbar_demux_035:sink_endofpacket
	wire         id_router_035_src_valid;                                                                           // id_router_035:src_valid -> rsp_xbar_demux_035:sink_valid
	wire         id_router_035_src_startofpacket;                                                                   // id_router_035:src_startofpacket -> rsp_xbar_demux_035:sink_startofpacket
	wire  [98:0] id_router_035_src_data;                                                                            // id_router_035:src_data -> rsp_xbar_demux_035:sink_data
	wire  [36:0] id_router_035_src_channel;                                                                         // id_router_035:src_channel -> rsp_xbar_demux_035:sink_channel
	wire         id_router_035_src_ready;                                                                           // rsp_xbar_demux_035:sink_ready -> id_router_035:src_ready
	wire         cmd_xbar_demux_001_src36_ready;                                                                    // switch8_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src36_ready
	wire         id_router_036_src_endofpacket;                                                                     // id_router_036:src_endofpacket -> rsp_xbar_demux_036:sink_endofpacket
	wire         id_router_036_src_valid;                                                                           // id_router_036:src_valid -> rsp_xbar_demux_036:sink_valid
	wire         id_router_036_src_startofpacket;                                                                   // id_router_036:src_startofpacket -> rsp_xbar_demux_036:sink_startofpacket
	wire  [98:0] id_router_036_src_data;                                                                            // id_router_036:src_data -> rsp_xbar_demux_036:sink_data
	wire  [36:0] id_router_036_src_channel;                                                                         // id_router_036:src_channel -> rsp_xbar_demux_036:sink_channel
	wire         id_router_036_src_ready;                                                                           // rsp_xbar_demux_036:sink_ready -> id_router_036:src_ready
	wire         crosser_out_endofpacket;                                                                           // crosser:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_out_valid;                                                                                 // crosser:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_out_startofpacket;                                                                         // crosser:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] crosser_out_data;                                                                                  // crosser:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] crosser_out_channel;                                                                               // crosser:out_channel -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src25_endofpacket;                                                              // cmd_xbar_demux_001:src25_endofpacket -> crosser:in_endofpacket
	wire         cmd_xbar_demux_001_src25_valid;                                                                    // cmd_xbar_demux_001:src25_valid -> crosser:in_valid
	wire         cmd_xbar_demux_001_src25_startofpacket;                                                            // cmd_xbar_demux_001:src25_startofpacket -> crosser:in_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src25_data;                                                                     // cmd_xbar_demux_001:src25_data -> crosser:in_data
	wire  [36:0] cmd_xbar_demux_001_src25_channel;                                                                  // cmd_xbar_demux_001:src25_channel -> crosser:in_channel
	wire         cmd_xbar_demux_001_src25_ready;                                                                    // crosser:in_ready -> cmd_xbar_demux_001:src25_ready
	wire         crosser_001_out_endofpacket;                                                                       // crosser_001:out_endofpacket -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_001_out_valid;                                                                             // crosser_001:out_valid -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_001_out_startofpacket;                                                                     // crosser_001:out_startofpacket -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [98:0] crosser_001_out_data;                                                                              // crosser_001:out_data -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [36:0] crosser_001_out_channel;                                                                           // crosser_001:out_channel -> clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src32_endofpacket;                                                              // cmd_xbar_demux_001:src32_endofpacket -> crosser_001:in_endofpacket
	wire         cmd_xbar_demux_001_src32_valid;                                                                    // cmd_xbar_demux_001:src32_valid -> crosser_001:in_valid
	wire         cmd_xbar_demux_001_src32_startofpacket;                                                            // cmd_xbar_demux_001:src32_startofpacket -> crosser_001:in_startofpacket
	wire  [98:0] cmd_xbar_demux_001_src32_data;                                                                     // cmd_xbar_demux_001:src32_data -> crosser_001:in_data
	wire  [36:0] cmd_xbar_demux_001_src32_channel;                                                                  // cmd_xbar_demux_001:src32_channel -> crosser_001:in_channel
	wire         cmd_xbar_demux_001_src32_ready;                                                                    // crosser_001:in_ready -> cmd_xbar_demux_001:src32_ready
	wire         crosser_002_out_endofpacket;                                                                       // crosser_002:out_endofpacket -> rsp_xbar_mux_001:sink25_endofpacket
	wire         crosser_002_out_valid;                                                                             // crosser_002:out_valid -> rsp_xbar_mux_001:sink25_valid
	wire         crosser_002_out_startofpacket;                                                                     // crosser_002:out_startofpacket -> rsp_xbar_mux_001:sink25_startofpacket
	wire  [98:0] crosser_002_out_data;                                                                              // crosser_002:out_data -> rsp_xbar_mux_001:sink25_data
	wire  [36:0] crosser_002_out_channel;                                                                           // crosser_002:out_channel -> rsp_xbar_mux_001:sink25_channel
	wire         crosser_002_out_ready;                                                                             // rsp_xbar_mux_001:sink25_ready -> crosser_002:out_ready
	wire         rsp_xbar_demux_025_src0_endofpacket;                                                               // rsp_xbar_demux_025:src0_endofpacket -> crosser_002:in_endofpacket
	wire         rsp_xbar_demux_025_src0_valid;                                                                     // rsp_xbar_demux_025:src0_valid -> crosser_002:in_valid
	wire         rsp_xbar_demux_025_src0_startofpacket;                                                             // rsp_xbar_demux_025:src0_startofpacket -> crosser_002:in_startofpacket
	wire  [98:0] rsp_xbar_demux_025_src0_data;                                                                      // rsp_xbar_demux_025:src0_data -> crosser_002:in_data
	wire  [36:0] rsp_xbar_demux_025_src0_channel;                                                                   // rsp_xbar_demux_025:src0_channel -> crosser_002:in_channel
	wire         rsp_xbar_demux_025_src0_ready;                                                                     // crosser_002:in_ready -> rsp_xbar_demux_025:src0_ready
	wire         crosser_003_out_endofpacket;                                                                       // crosser_003:out_endofpacket -> rsp_xbar_mux_001:sink32_endofpacket
	wire         crosser_003_out_valid;                                                                             // crosser_003:out_valid -> rsp_xbar_mux_001:sink32_valid
	wire         crosser_003_out_startofpacket;                                                                     // crosser_003:out_startofpacket -> rsp_xbar_mux_001:sink32_startofpacket
	wire  [98:0] crosser_003_out_data;                                                                              // crosser_003:out_data -> rsp_xbar_mux_001:sink32_data
	wire  [36:0] crosser_003_out_channel;                                                                           // crosser_003:out_channel -> rsp_xbar_mux_001:sink32_channel
	wire         crosser_003_out_ready;                                                                             // rsp_xbar_mux_001:sink32_ready -> crosser_003:out_ready
	wire         rsp_xbar_demux_032_src0_endofpacket;                                                               // rsp_xbar_demux_032:src0_endofpacket -> crosser_003:in_endofpacket
	wire         rsp_xbar_demux_032_src0_valid;                                                                     // rsp_xbar_demux_032:src0_valid -> crosser_003:in_valid
	wire         rsp_xbar_demux_032_src0_startofpacket;                                                             // rsp_xbar_demux_032:src0_startofpacket -> crosser_003:in_startofpacket
	wire  [98:0] rsp_xbar_demux_032_src0_data;                                                                      // rsp_xbar_demux_032:src0_data -> crosser_003:in_data
	wire  [36:0] rsp_xbar_demux_032_src0_channel;                                                                   // rsp_xbar_demux_032:src0_channel -> crosser_003:in_channel
	wire         rsp_xbar_demux_032_src0_ready;                                                                     // crosser_003:in_ready -> rsp_xbar_demux_032:src0_ready
	wire  [36:0] limiter_cmd_valid_data;                                                                            // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire  [36:0] limiter_001_cmd_valid_data;                                                                        // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                          // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                          // uart:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                          // bclk_out:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                          // lrcin:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                                          // key1:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                                          // key2:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                                                          // key3:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                                                          // switch0:irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                                                          // key0:irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                                                                          // switch1:irq -> irq_mapper:receiver9_irq
	wire         irq_mapper_receiver10_irq;                                                                         // switch2:irq -> irq_mapper:receiver10_irq
	wire         irq_mapper_receiver11_irq;                                                                         // switch3:irq -> irq_mapper:receiver11_irq
	wire         irq_mapper_receiver12_irq;                                                                         // switch4:irq -> irq_mapper:receiver12_irq
	wire         irq_mapper_receiver13_irq;                                                                         // leftready:irq -> irq_mapper:receiver13_irq
	wire         irq_mapper_receiver14_irq;                                                                         // rightready:irq -> irq_mapper:receiver14_irq
	wire         irq_mapper_receiver15_irq;                                                                         // bclk_in:irq -> irq_mapper:receiver15_irq
	wire         irq_mapper_receiver16_irq;                                                                         // lrcout:irq -> irq_mapper:receiver16_irq
	wire         irq_mapper_receiver17_irq;                                                                         // switch5:irq -> irq_mapper:receiver17_irq
	wire         irq_mapper_receiver18_irq;                                                                         // switch6:irq -> irq_mapper:receiver18_irq
	wire         irq_mapper_receiver19_irq;                                                                         // switch7:irq -> irq_mapper:receiver19_irq
	wire         irq_mapper_receiver20_irq;                                                                         // switch8:irq -> irq_mapper:receiver20_irq
	wire  [31:0] nios2_qsys_d_irq_irq;                                                                              // irq_mapper:sender_irq -> nios2_qsys:d_irq

	de2i_150_nios2_qsys nios2_qsys (
		.clk                                   (altpll_0_c0_clk),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                         //                   reset_n.reset_n
		.d_address                             (nios2_qsys_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                                        //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                         // custom_instruction_master.readra
	);

	de2i_150_uart uart (
		.clk           (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address       (uart_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                     //                    .dataavailable
		.readyfordata  (),                                                     //                    .readyfordata
		.rxd           (uart_rxd),                                             // external_connection.export
		.txd           (uart_txd),                                             //                    .export
		.irq           (irq_mapper_receiver1_irq)                              //                 irq.irq
	);

	de2i_150_jtag_uart jtag_uart (
		.clk            (altpll_0_c0_clk),                                                        //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	de2i_150_sysid_qsys sysid_qsys (
		.clock    (altpll_0_c0_clk),                                                  //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                  //         reset.reset_n
		.readdata (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	de2i_150_led led (
		.clk        (altpll_0_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_export)                                        // external_connection.export
	);

	de2i_150_switch0 switch0 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch0_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver7_irq)                              //                 irq.irq
	);

	de2i_150_key0 key0 (
		.clk        (altpll_0_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (key0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~key0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (key0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (key0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (key0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key0_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver8_irq)                           //                 irq.irq
	);

	de2i_150_onchip_memory2 onchip_memory2 (
		.clk        (altpll_0_c0_clk),                                             //   clk1.clk
		.address    (onchip_memory2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                           //       .reset_req
	);

	de2i_150_adc adc (
		.clk      (altpll_0_c0_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (adc_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (adc_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (adc_export)                                      // external_connection.export
	);

	de2i_150_cs cs (
		.clk        (altpll_0_c0_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (cs_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~cs_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (cs_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (cs_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (cs_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (cs_export)                                        // external_connection.export
	);

	de2i_150_cs sclk (
		.clk        (altpll_0_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (sclk_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sclk_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sclk_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sclk_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sclk_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (sclk_export)                                        // external_connection.export
	);

	de2i_150_cs sdin (
		.clk        (altpll_0_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (sdin_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~sdin_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (sdin_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (sdin_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (sdin_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (sdin_export)                                        // external_connection.export
	);

	de2i_150_cs din (
		.clk        (altpll_0_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (din_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~din_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (din_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (din_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (din_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (din_export)                                        // external_connection.export
	);

	de2i_150_key0 bclk_in (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (bclk_in_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~bclk_in_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (bclk_in_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (bclk_in_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (bclk_in_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (bclk_in_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver15_irq)                             //                 irq.irq
	);

	de2i_150_switch0 lrcout (
		.clk        (altpll_0_c0_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (lrcout_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lrcout_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lrcout_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lrcout_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lrcout_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (lrcout_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver16_irq)                            //                 irq.irq
	);

	de2i_150_dout dout (
		.clk      (altpll_0_c0_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (dout_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (dout_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (dout_export)                                      // external_connection.export
	);

	de2i_150_key0 bclk_out (
		.clk        (altpll_0_c0_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (bclk_out_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~bclk_out_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (bclk_out_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (bclk_out_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (bclk_out_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (bclk_out_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                               //                 irq.irq
	);

	de2i_150_switch0 lrcin (
		.clk        (altpll_0_c0_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (lrcin_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lrcin_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lrcin_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lrcin_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lrcin_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (lrcin_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                            //                 irq.irq
	);

	de2i_150_key0 key1 (
		.clk        (altpll_0_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (key1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~key1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (key1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (key1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (key1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key1_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                           //                 irq.irq
	);

	de2i_150_key0 key2 (
		.clk        (altpll_0_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (key2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~key2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (key2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (key2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (key2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key2_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                           //                 irq.irq
	);

	de2i_150_key0 key3 (
		.clk        (altpll_0_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (key3_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~key3_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (key3_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (key3_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (key3_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key3_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver6_irq)                           //                 irq.irq
	);

	de2i_150_switch0 switch1 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch1_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver9_irq)                              //                 irq.irq
	);

	de2i_150_switch0 switch2 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch2_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver10_irq)                             //                 irq.irq
	);

	de2i_150_switch0 switch3 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch3_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch3_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch3_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch3_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch3_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch3_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver11_irq)                             //                 irq.irq
	);

	de2i_150_switch0 switch4 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch4_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch4_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch4_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch4_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch4_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch4_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver12_irq)                             //                 irq.irq
	);

	de2i_150_altpll_0 altpll_0 (
		.clk       (clk_clk),                                                     //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),                          // inclk_interface_reset.reset
		.read      (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (altpll_0_c0_clk),                                             //                    c0.clk
		.areset    (),                                                            //        areset_conduit.export
		.locked    (),                                                            //        locked_conduit.export
		.phasedone ()                                                             //     phasedone_conduit.export
	);

	de2i_150_leftdata leftdata (
		.clk      (altpll_0_c0_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address  (leftdata_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (leftdata_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (leftdata_export)                                      // external_connection.export
	);

	de2i_150_leftdata rightdata (
		.clk      (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address  (rightdata_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (rightdata_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (rightdata_export)                                      // external_connection.export
	);

	de2i_150_key0 leftready (
		.clk        (altpll_0_c0_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (leftready_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~leftready_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (leftready_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (leftready_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (leftready_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (leftready_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver13_irq)                               //                 irq.irq
	);

	de2i_150_key0 rightready (
		.clk        (altpll_0_c0_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (rightready_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~rightready_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (rightready_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (rightready_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (rightready_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (rightready_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver14_irq)                                //                 irq.irq
	);

	de2i_150_leftsenddata leftsenddata (
		.clk        (altpll_0_c0_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           //               reset.reset_n
		.address    (leftsenddata_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~leftsenddata_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (leftsenddata_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (leftsenddata_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (leftsenddata_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (leftsenddata_export)                                        // external_connection.export
	);

	de2i_150_leftsenddata rightsenddata (
		.clk        (altpll_0_c0_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //               reset.reset_n
		.address    (rightsenddata_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~rightsenddata_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (rightsenddata_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (rightsenddata_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (rightsenddata_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (rightsenddata_export)                                        // external_connection.export
	);

	de2i_150_clk_12mhz clk_12mhz (
		.clk       (clk_clk),                                                      //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),                           // inclk_interface_reset.reset
		.read      (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (clk_12mhz_c0_clk),                                             //                    c0.clk
		.areset    (),                                                             //        areset_conduit.export
		.locked    (),                                                             //        locked_conduit.export
		.phasedone ()                                                              //     phasedone_conduit.export
	);

	de2i_150_switch0 switch5 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch5_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch5_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch5_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch5_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch5_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch5_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver17_irq)                             //                 irq.irq
	);

	de2i_150_switch6 switch6 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch6_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch6_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch6_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch6_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch6_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch6_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver18_irq)                             //                 irq.irq
	);

	de2i_150_switch0 switch7 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch7_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch7_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch7_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch7_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch7_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch7_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver19_irq)                             //                 irq.irq
	);

	de2i_150_switch0 switch8 (
		.clk        (altpll_0_c0_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (switch8_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~switch8_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (switch8_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (switch8_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (switch8_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (switch8_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver20_irq)                             //                 irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (20),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (20),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_instruction_master_translator (
		.clk                      (altpll_0_c0_clk),                                                                  //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_qsys_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                             //               (terminated)
		.av_byteenable            (4'b1111),                                                                          //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                             //               (terminated)
		.av_begintransfer         (1'b0),                                                                             //               (terminated)
		.av_chipselect            (1'b0),                                                                             //               (terminated)
		.av_write                 (1'b0),                                                                             //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                             //               (terminated)
		.av_lock                  (1'b0),                                                                             //               (terminated)
		.av_debugaccess           (1'b0),                                                                             //               (terminated)
		.uav_clken                (),                                                                                 //               (terminated)
		.av_clken                 (1'b1),                                                                             //               (terminated)
		.uav_response             (2'b00),                                                                            //               (terminated)
		.av_response              (),                                                                                 //               (terminated)
		.uav_writeresponserequest (),                                                                                 //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                             //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                             //               (terminated)
		.av_writeresponsevalid    ()                                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (20),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (20),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_data_master_translator (
		.clk                      (altpll_0_c0_clk),                                                           //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (nios2_qsys_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_qsys_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_qsys_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (nios2_qsys_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_jtag_debug_module_translator (
		.clk                      (altpll_0_c0_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                                        //              (terminated)
		.av_burstcount            (),                                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                        //              (terminated)
		.av_lock                  (),                                                                                        //              (terminated)
		.av_chipselect            (),                                                                                        //              (terminated)
		.av_clken                 (),                                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                        //              (terminated)
		.uav_response             (),                                                                                        //              (terminated)
		.av_response              (2'b00),                                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (16),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (uart_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_control_slave_translator (
		.clk                      (altpll_0_c0_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                                    //              (terminated)
		.av_read                  (),                                                                                    //              (terminated)
		.av_writedata             (),                                                                                    //              (terminated)
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch0_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key0_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (key0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (key0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (key0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (key0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (key0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) adc_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (adc_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (adc_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (adc_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (adc_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (adc_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (adc_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (adc_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (adc_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (adc_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (adc_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (adc_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (adc_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (adc_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                  //              (terminated)
		.av_read                  (),                                                                  //              (terminated)
		.av_writedata             (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_chipselect            (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cs_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                   //                    reset.reset
		.uav_address              (cs_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cs_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cs_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cs_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cs_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cs_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cs_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cs_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (cs_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cs_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (cs_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                 //              (terminated)
		.av_begintransfer         (),                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                 //              (terminated)
		.av_burstcount            (),                                                                 //              (terminated)
		.av_byteenable            (),                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                             //              (terminated)
		.av_writebyteenable       (),                                                                 //              (terminated)
		.av_lock                  (),                                                                 //              (terminated)
		.av_clken                 (),                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                             //              (terminated)
		.av_debugaccess           (),                                                                 //              (terminated)
		.av_outputenable          (),                                                                 //              (terminated)
		.uav_response             (),                                                                 //              (terminated)
		.av_response              (2'b00),                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sclk_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (sclk_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sclk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sclk_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sclk_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sclk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sclk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sclk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sclk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sclk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sclk_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sclk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sclk_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sclk_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (sclk_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sclk_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sclk_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdin_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (sdin_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdin_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdin_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdin_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdin_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdin_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdin_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdin_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (sdin_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdin_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sdin_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) din_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (din_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (din_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (din_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (din_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (din_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (din_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (din_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (din_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (din_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (din_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (din_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (din_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (din_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (din_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (din_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (din_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) bclk_in_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (bclk_in_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (bclk_in_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (bclk_in_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (bclk_in_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (bclk_in_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lrcout_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lrcout_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lrcout_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lrcout_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lrcout_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lrcout_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dout_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (dout_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dout_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dout_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dout_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dout_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dout_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dout_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (dout_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                   //              (terminated)
		.av_read                  (),                                                                   //              (terminated)
		.av_writedata             (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_chipselect            (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) bclk_out_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (bclk_out_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (bclk_out_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (bclk_out_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (bclk_out_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (bclk_out_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lrcin_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lrcin_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lrcin_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lrcin_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lrcin_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lrcin_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key1_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (key1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (key1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (key1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (key1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (key1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key2_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (key2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (key2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (key2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (key2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (key2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key3_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (key3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (key3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (key3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (key3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (key3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch1_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch2_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch3_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch4_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altpll_0_pll_slave_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leftdata_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (leftdata_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (leftdata_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rightdata_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (rightdata_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (rightdata_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                        //              (terminated)
		.av_read                  (),                                                                        //              (terminated)
		.av_writedata             (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_chipselect            (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leftready_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (leftready_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (leftready_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (leftready_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (leftready_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (leftready_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (leftready_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (leftready_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (leftready_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (leftready_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (leftready_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (leftready_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (leftready_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (leftready_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (leftready_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (leftready_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (leftready_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rightready_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address              (rightready_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (rightready_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (rightready_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (rightready_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (rightready_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (rightready_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (rightready_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (rightready_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (rightready_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (rightready_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (rightready_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (rightready_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (rightready_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (rightready_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (rightready_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (rightready_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leftsenddata_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address              (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (leftsenddata_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (leftsenddata_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (leftsenddata_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (leftsenddata_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (leftsenddata_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rightsenddata_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address              (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (rightsenddata_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (rightsenddata_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (rightsenddata_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (rightsenddata_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (rightsenddata_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) clk_12mhz_pll_slave_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (clk_12mhz_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch5_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch6_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch6_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch6_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch6_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch6_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch6_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch6_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch6_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch6_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch6_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch7_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch7_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch7_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch7_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch7_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch7_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch7_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch7_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch7_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch7_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch8_s1_translator (
		.clk                      (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (switch8_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch8_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch8_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch8_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch8_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch8_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch8_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch8_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch8_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch8_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch8_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch8_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (switch8_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (switch8_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (switch8_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (switch8_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_BEGIN_BURST           (75),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.PKT_BURST_TYPE_H          (72),
		.PKT_BURST_TYPE_L          (71),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_TRANS_EXCLUSIVE       (61),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_THREAD_ID_H           (89),
		.PKT_THREAD_ID_L           (89),
		.PKT_CACHE_H               (96),
		.PKT_CACHE_L               (93),
		.PKT_DATA_SIDEBAND_H       (74),
		.PKT_DATA_SIDEBAND_L       (74),
		.PKT_QOS_H                 (76),
		.PKT_QOS_L                 (76),
		.PKT_ADDR_SIDEBAND_H       (73),
		.PKT_ADDR_SIDEBAND_L       (73),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (37),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                           //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.av_address              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                                     //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                                      //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                                   //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                             //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                               //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                                     //          .ready
		.av_response             (),                                                                                          // (terminated)
		.av_writeresponserequest (1'b0),                                                                                      // (terminated)
		.av_writeresponsevalid   ()                                                                                           // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_BEGIN_BURST           (75),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.PKT_BURST_TYPE_H          (72),
		.PKT_BURST_TYPE_L          (71),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_TRANS_EXCLUSIVE       (61),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_THREAD_ID_H           (89),
		.PKT_THREAD_ID_L           (89),
		.PKT_CACHE_H               (96),
		.PKT_CACHE_L               (93),
		.PKT_DATA_SIDEBAND_H       (74),
		.PKT_DATA_SIDEBAND_L       (74),
		.PKT_QOS_H                 (76),
		.PKT_QOS_L                 (76),
		.PKT_ADDR_SIDEBAND_H       (73),
		.PKT_ADDR_SIDEBAND_L       (73),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (37),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (nios2_qsys_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                          //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                           //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                          //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                          //                .channel
		.rf_sink_ready           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                           //                .channel
		.rf_sink_ready           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (uart_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                              //                .channel
		.rf_sink_ready           (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                               //                .channel
		.rf_sink_ready           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                             //                .channel
		.rf_sink_ready           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                 //                .channel
		.rf_sink_ready           (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (key0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                              //                .channel
		.rf_sink_ready           (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) adc_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (adc_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (adc_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (adc_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (adc_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (adc_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (adc_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (adc_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (adc_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (adc_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (adc_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (adc_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (adc_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (adc_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (adc_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (adc_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (adc_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                             //                .channel
		.rf_sink_ready           (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (adc_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (adc_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (adc_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cs_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (cs_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cs_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cs_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cs_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cs_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cs_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cs_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cs_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cs_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                            //                .channel
		.rf_sink_ready           (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.in_data           (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sclk_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (sclk_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sclk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sclk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sclk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sclk_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sclk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sclk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sclk_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sclk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sclk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sclk_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sclk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sclk_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sclk_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sclk_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sclk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                             //                .channel
		.rf_sink_ready           (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sclk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdin_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (sdin_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdin_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdin_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdin_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdin_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdin_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdin_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdin_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdin_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                             //                .channel
		.rf_sink_ready           (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) din_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (din_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (din_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (din_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (din_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (din_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (din_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (din_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (din_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (din_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (din_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (din_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (din_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (din_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (din_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (din_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (din_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                              //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                            //                .channel
		.rf_sink_ready           (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (din_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (din_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (din_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (din_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (din_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (din_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (din_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (din_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (din_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (din_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (din_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (din_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) bclk_in_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (bclk_in_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                //                .channel
		.rf_sink_ready           (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (bclk_in_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (bclk_in_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (bclk_in_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lrcout_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lrcout_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                               //                .channel
		.rf_sink_ready           (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lrcout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lrcout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lrcout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dout_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (dout_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dout_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dout_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dout_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dout_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dout_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dout_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dout_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dout_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dout_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dout_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dout_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dout_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dout_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                             //                .channel
		.rf_sink_ready           (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dout_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dout_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dout_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) bclk_out_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (bclk_out_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                 //                .channel
		.rf_sink_ready           (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (bclk_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (bclk_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (bclk_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lrcin_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lrcin_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                              //                .channel
		.rf_sink_ready           (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lrcin_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lrcin_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lrcin_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (key1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                             //                .channel
		.rf_sink_ready           (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (key2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src19_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src19_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src19_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src19_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src19_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src19_channel),                                             //                .channel
		.rf_sink_ready           (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (key3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src20_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src20_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src20_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src20_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src20_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src20_channel),                                             //                .channel
		.rf_sink_ready           (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src21_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src21_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src21_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src21_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src21_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src21_channel),                                                //                .channel
		.rf_sink_ready           (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src22_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src22_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src22_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src22_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src22_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src22_channel),                                                //                .channel
		.rf_sink_ready           (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src23_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src23_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src23_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src23_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src23_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src23_channel),                                                //                .channel
		.rf_sink_ready           (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src24_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src24_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src24_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src24_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src24_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src24_channel),                                                //                .channel
		.rf_sink_ready           (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                       //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                       //                .valid
		.cp_data                 (crosser_out_data),                                                                        //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                     //                .channel
		.rf_sink_ready           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) leftdata_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leftdata_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src26_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src26_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src26_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src26_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src26_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src26_channel),                                                 //                .channel
		.rf_sink_ready           (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leftdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leftdata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leftdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rightdata_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rightdata_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src27_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src27_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src27_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src27_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src27_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src27_channel),                                                  //                .channel
		.rf_sink_ready           (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rightdata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rightdata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rightdata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) leftready_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (leftready_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leftready_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leftready_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leftready_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leftready_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leftready_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leftready_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leftready_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leftready_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leftready_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leftready_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leftready_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leftready_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leftready_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leftready_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leftready_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src28_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src28_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src28_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src28_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src28_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src28_channel),                                                  //                .channel
		.rf_sink_ready           (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leftready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leftready_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leftready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rightready_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (rightready_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rightready_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rightready_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rightready_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rightready_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rightready_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rightready_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rightready_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rightready_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rightready_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rightready_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rightready_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rightready_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rightready_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rightready_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rightready_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src29_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src29_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src29_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src29_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src29_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src29_channel),                                                   //                .channel
		.rf_sink_ready           (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rightready_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rightready_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rightready_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) leftsenddata_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leftsenddata_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src30_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src30_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src30_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src30_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src30_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src30_channel),                                                     //                .channel
		.rf_sink_ready           (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rightsenddata_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rightsenddata_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src31_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src31_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src31_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src31_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src31_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src31_channel),                                                      //                .channel
		.rf_sink_ready           (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_001_out_ready),                                                                    //              cp.ready
		.cp_valid                (crosser_001_out_valid),                                                                    //                .valid
		.cp_data                 (crosser_001_out_data),                                                                     //                .data
		.cp_startofpacket        (crosser_001_out_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (crosser_001_out_endofpacket),                                                              //                .endofpacket
		.cp_channel              (crosser_001_out_channel),                                                                  //                .channel
		.rf_sink_ready           (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_startofpacket  (1'b0),                                                                               // (terminated)
		.in_endofpacket    (1'b0),                                                                               // (terminated)
		.out_startofpacket (),                                                                                   // (terminated)
		.out_endofpacket   (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src33_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src33_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src33_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src33_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src33_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src33_channel),                                                //                .channel
		.rf_sink_ready           (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch6_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch6_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch6_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch6_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch6_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch6_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch6_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch6_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src34_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src34_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src34_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src34_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src34_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src34_channel),                                                //                .channel
		.rf_sink_ready           (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch7_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch7_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch7_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch7_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch7_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch7_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch7_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch7_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src35_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src35_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src35_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src35_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src35_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src35_channel),                                                //                .channel
		.rf_sink_ready           (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (77),
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (67),
		.PKT_BURSTWRAP_L           (65),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (90),
		.PKT_RESPONSE_STATUS_H     (98),
		.PKT_RESPONSE_STATUS_L     (97),
		.PKT_BURST_SIZE_H          (70),
		.PKT_BURST_SIZE_L          (68),
		.ST_CHANNEL_W              (37),
		.ST_DATA_W                 (99),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch8_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (switch8_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch8_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch8_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch8_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch8_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch8_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch8_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch8_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch8_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch8_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch8_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch8_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch8_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch8_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch8_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch8_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src36_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src36_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src36_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src36_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src36_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src36_channel),                                                //                .channel
		.rf_sink_ready           (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch8_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (100),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch8_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch8_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	de2i_150_addr_router addr_router (
		.sink_ready         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                     //       src.ready
		.src_valid          (addr_router_src_valid),                                                                     //          .valid
		.src_data           (addr_router_src_data),                                                                      //          .data
		.src_channel        (addr_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                //          .endofpacket
	);

	de2i_150_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                          //          .valid
		.src_data           (addr_router_001_src_data),                                                           //          .data
		.src_channel        (addr_router_001_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                     //          .endofpacket
	);

	de2i_150_id_router id_router (
		.sink_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_src_valid),                                                                     //          .valid
		.src_data           (id_router_src_data),                                                                      //          .data
		.src_channel        (id_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                //          .endofpacket
	);

	de2i_150_id_router id_router_001 (
		.sink_ready         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                      //       src.ready
		.src_valid          (id_router_001_src_valid),                                                      //          .valid
		.src_data           (id_router_001_src_data),                                                       //          .data
		.src_channel        (id_router_001_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                 //          .endofpacket
	);

	de2i_150_id_router_002 id_router_002 (
		.sink_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                            //       src.ready
		.src_valid          (id_router_002_src_valid),                                            //          .valid
		.src_data           (id_router_002_src_data),                                             //          .data
		.src_channel        (id_router_002_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                       //          .endofpacket
	);

	de2i_150_id_router_002 id_router_003 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                //          .valid
		.src_data           (id_router_003_src_data),                                                                 //          .data
		.src_channel        (id_router_003_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                           //          .endofpacket
	);

	de2i_150_id_router_002 id_router_004 (
		.sink_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                             //       src.ready
		.src_valid          (id_router_004_src_valid),                                                             //          .valid
		.src_data           (id_router_004_src_data),                                                              //          .data
		.src_channel        (id_router_004_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                        //          .endofpacket
	);

	de2i_150_id_router_002 id_router_005 (
		.sink_ready         (led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                           //       src.ready
		.src_valid          (id_router_005_src_valid),                                           //          .valid
		.src_data           (id_router_005_src_data),                                            //          .data
		.src_channel        (id_router_005_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                      //          .endofpacket
	);

	de2i_150_id_router_002 id_router_006 (
		.sink_ready         (switch0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                               //       src.ready
		.src_valid          (id_router_006_src_valid),                                               //          .valid
		.src_data           (id_router_006_src_data),                                                //          .data
		.src_channel        (id_router_006_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_007 (
		.sink_ready         (key0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                            //       src.ready
		.src_valid          (id_router_007_src_valid),                                            //          .valid
		.src_data           (id_router_007_src_data),                                             //          .data
		.src_channel        (id_router_007_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                       //          .endofpacket
	);

	de2i_150_id_router_002 id_router_008 (
		.sink_ready         (adc_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (adc_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (adc_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (adc_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (adc_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                           //       src.ready
		.src_valid          (id_router_008_src_valid),                                           //          .valid
		.src_data           (id_router_008_src_data),                                            //          .data
		.src_channel        (id_router_008_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                      //          .endofpacket
	);

	de2i_150_id_router_002 id_router_009 (
		.sink_ready         (cs_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cs_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cs_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                          //       src.ready
		.src_valid          (id_router_009_src_valid),                                          //          .valid
		.src_data           (id_router_009_src_data),                                           //          .data
		.src_channel        (id_router_009_src_channel),                                        //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                  //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                     //          .endofpacket
	);

	de2i_150_id_router_002 id_router_010 (
		.sink_ready         (sclk_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sclk_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sclk_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sclk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sclk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                            //       src.ready
		.src_valid          (id_router_010_src_valid),                                            //          .valid
		.src_data           (id_router_010_src_data),                                             //          .data
		.src_channel        (id_router_010_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                       //          .endofpacket
	);

	de2i_150_id_router_002 id_router_011 (
		.sink_ready         (sdin_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdin_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdin_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                            //       src.ready
		.src_valid          (id_router_011_src_valid),                                            //          .valid
		.src_data           (id_router_011_src_data),                                             //          .data
		.src_channel        (id_router_011_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                       //          .endofpacket
	);

	de2i_150_id_router_002 id_router_012 (
		.sink_ready         (din_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (din_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (din_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (din_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (din_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                           //       src.ready
		.src_valid          (id_router_012_src_valid),                                           //          .valid
		.src_data           (id_router_012_src_data),                                            //          .data
		.src_channel        (id_router_012_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                      //          .endofpacket
	);

	de2i_150_id_router_002 id_router_013 (
		.sink_ready         (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (bclk_in_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                               //       src.ready
		.src_valid          (id_router_013_src_valid),                                               //          .valid
		.src_data           (id_router_013_src_data),                                                //          .data
		.src_channel        (id_router_013_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_014 (
		.sink_ready         (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lrcout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                              //       src.ready
		.src_valid          (id_router_014_src_valid),                                              //          .valid
		.src_data           (id_router_014_src_data),                                               //          .data
		.src_channel        (id_router_014_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                         //          .endofpacket
	);

	de2i_150_id_router_002 id_router_015 (
		.sink_ready         (dout_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dout_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dout_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dout_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dout_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                            //       src.ready
		.src_valid          (id_router_015_src_valid),                                            //          .valid
		.src_data           (id_router_015_src_data),                                             //          .data
		.src_channel        (id_router_015_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                       //          .endofpacket
	);

	de2i_150_id_router_002 id_router_016 (
		.sink_ready         (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (bclk_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                //       src.ready
		.src_valid          (id_router_016_src_valid),                                                //          .valid
		.src_data           (id_router_016_src_data),                                                 //          .data
		.src_channel        (id_router_016_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                           //          .endofpacket
	);

	de2i_150_id_router_002 id_router_017 (
		.sink_ready         (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lrcin_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                             //       src.ready
		.src_valid          (id_router_017_src_valid),                                             //          .valid
		.src_data           (id_router_017_src_data),                                              //          .data
		.src_channel        (id_router_017_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                        //          .endofpacket
	);

	de2i_150_id_router_002 id_router_018 (
		.sink_ready         (key1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                            //       src.ready
		.src_valid          (id_router_018_src_valid),                                            //          .valid
		.src_data           (id_router_018_src_data),                                             //          .data
		.src_channel        (id_router_018_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                       //          .endofpacket
	);

	de2i_150_id_router_002 id_router_019 (
		.sink_ready         (key2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                            //       src.ready
		.src_valid          (id_router_019_src_valid),                                            //          .valid
		.src_data           (id_router_019_src_data),                                             //          .data
		.src_channel        (id_router_019_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                       //          .endofpacket
	);

	de2i_150_id_router_002 id_router_020 (
		.sink_ready         (key3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                            //       src.ready
		.src_valid          (id_router_020_src_valid),                                            //          .valid
		.src_data           (id_router_020_src_data),                                             //          .data
		.src_channel        (id_router_020_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                       //          .endofpacket
	);

	de2i_150_id_router_002 id_router_021 (
		.sink_ready         (switch1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                               //       src.ready
		.src_valid          (id_router_021_src_valid),                                               //          .valid
		.src_data           (id_router_021_src_data),                                                //          .data
		.src_channel        (id_router_021_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_022 (
		.sink_ready         (switch2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                               //       src.ready
		.src_valid          (id_router_022_src_valid),                                               //          .valid
		.src_data           (id_router_022_src_data),                                                //          .data
		.src_channel        (id_router_022_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_023 (
		.sink_ready         (switch3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                               //       src.ready
		.src_valid          (id_router_023_src_valid),                                               //          .valid
		.src_data           (id_router_023_src_data),                                                //          .data
		.src_channel        (id_router_023_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_024 (
		.sink_ready         (switch4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                               //       src.ready
		.src_valid          (id_router_024_src_valid),                                               //          .valid
		.src_data           (id_router_024_src_data),                                                //          .data
		.src_channel        (id_router_024_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_025 (
		.sink_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                       //       src.ready
		.src_valid          (id_router_025_src_valid),                                                       //          .valid
		.src_data           (id_router_025_src_data),                                                        //          .data
		.src_channel        (id_router_025_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                                  //          .endofpacket
	);

	de2i_150_id_router_002 id_router_026 (
		.sink_ready         (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leftdata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                //       src.ready
		.src_valid          (id_router_026_src_valid),                                                //          .valid
		.src_data           (id_router_026_src_data),                                                 //          .data
		.src_channel        (id_router_026_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                           //          .endofpacket
	);

	de2i_150_id_router_002 id_router_027 (
		.sink_ready         (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rightdata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                 //       src.ready
		.src_valid          (id_router_027_src_valid),                                                 //          .valid
		.src_data           (id_router_027_src_data),                                                  //          .data
		.src_channel        (id_router_027_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                            //          .endofpacket
	);

	de2i_150_id_router_002 id_router_028 (
		.sink_ready         (leftready_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leftready_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leftready_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leftready_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leftready_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                                 //       src.ready
		.src_valid          (id_router_028_src_valid),                                                 //          .valid
		.src_data           (id_router_028_src_data),                                                  //          .data
		.src_channel        (id_router_028_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                            //          .endofpacket
	);

	de2i_150_id_router_002 id_router_029 (
		.sink_ready         (rightready_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rightready_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rightready_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rightready_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rightready_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                  //       src.ready
		.src_valid          (id_router_029_src_valid),                                                  //          .valid
		.src_data           (id_router_029_src_data),                                                   //          .data
		.src_channel        (id_router_029_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                             //          .endofpacket
	);

	de2i_150_id_router_002 id_router_030 (
		.sink_ready         (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leftsenddata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                                    //       src.ready
		.src_valid          (id_router_030_src_valid),                                                    //          .valid
		.src_data           (id_router_030_src_data),                                                     //          .data
		.src_channel        (id_router_030_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                               //          .endofpacket
	);

	de2i_150_id_router_002 id_router_031 (
		.sink_ready         (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rightsenddata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                                     //       src.ready
		.src_valid          (id_router_031_src_valid),                                                     //          .valid
		.src_data           (id_router_031_src_data),                                                      //          .data
		.src_channel        (id_router_031_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                                //          .endofpacket
	);

	de2i_150_id_router_002 id_router_032 (
		.sink_ready         (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (clk_12mhz_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                                        //       src.ready
		.src_valid          (id_router_032_src_valid),                                                        //          .valid
		.src_data           (id_router_032_src_data),                                                         //          .data
		.src_channel        (id_router_032_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                                   //          .endofpacket
	);

	de2i_150_id_router_002 id_router_033 (
		.sink_ready         (switch5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_033_src_ready),                                               //       src.ready
		.src_valid          (id_router_033_src_valid),                                               //          .valid
		.src_data           (id_router_033_src_data),                                                //          .data
		.src_channel        (id_router_033_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_033_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_033_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_034 (
		.sink_ready         (switch6_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch6_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch6_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_034_src_ready),                                               //       src.ready
		.src_valid          (id_router_034_src_valid),                                               //          .valid
		.src_data           (id_router_034_src_data),                                                //          .data
		.src_channel        (id_router_034_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_034_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_034_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_035 (
		.sink_ready         (switch7_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch7_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch7_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_035_src_ready),                                               //       src.ready
		.src_valid          (id_router_035_src_valid),                                               //          .valid
		.src_data           (id_router_035_src_data),                                                //          .data
		.src_channel        (id_router_035_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_035_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_035_src_endofpacket)                                          //          .endofpacket
	);

	de2i_150_id_router_002 id_router_036 (
		.sink_ready         (switch8_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch8_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch8_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch8_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch8_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_036_src_ready),                                               //       src.ready
		.src_valid          (id_router_036_src_valid),                                               //          .valid
		.src_data           (id_router_036_src_data),                                                //          .data
		.src_channel        (id_router_036_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_036_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_036_src_endofpacket)                                          //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (37),
		.VALID_WIDTH               (37),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (altpll_0_c0_clk),                //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (88),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (99),
		.ST_CHANNEL_W              (37),
		.VALID_WIDTH               (37),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (64),
		.PKT_BYTE_CNT_L            (62),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (altpll_0_c0_clk),                    //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                           // reset_in0.reset
		.reset_in1  (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (altpll_0_c0_clk),                          //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_in2  (1'b0),                                     // (terminated)
		.reset_in3  (1'b0),                                     // (terminated)
		.reset_in4  (1'b0),                                     // (terminated)
		.reset_in5  (1'b0),                                     // (terminated)
		.reset_in6  (1'b0),                                     // (terminated)
		.reset_in7  (1'b0),                                     // (terminated)
		.reset_in8  (1'b0),                                     // (terminated)
		.reset_in9  (1'b0),                                     // (terminated)
		.reset_in10 (1'b0),                                     // (terminated)
		.reset_in11 (1'b0),                                     // (terminated)
		.reset_in12 (1'b0),                                     // (terminated)
		.reset_in13 (1'b0),                                     // (terminated)
		.reset_in14 (1'b0),                                     // (terminated)
		.reset_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	de2i_150_cmd_xbar_demux cmd_xbar_demux (
		.clk                (altpll_0_c0_clk),                   //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	de2i_150_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (altpll_0_c0_clk),                        //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //           .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //      src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //           .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //           .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //           .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //           .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //           .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //      src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //           .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //           .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //           .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //           .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //           .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //      src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //           .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //           .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //           .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //           .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //           .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //      src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //           .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //           .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //           .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //           .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket),   //           .endofpacket
		.src23_ready         (cmd_xbar_demux_001_src23_ready),         //      src23.ready
		.src23_valid         (cmd_xbar_demux_001_src23_valid),         //           .valid
		.src23_data          (cmd_xbar_demux_001_src23_data),          //           .data
		.src23_channel       (cmd_xbar_demux_001_src23_channel),       //           .channel
		.src23_startofpacket (cmd_xbar_demux_001_src23_startofpacket), //           .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_001_src23_endofpacket),   //           .endofpacket
		.src24_ready         (cmd_xbar_demux_001_src24_ready),         //      src24.ready
		.src24_valid         (cmd_xbar_demux_001_src24_valid),         //           .valid
		.src24_data          (cmd_xbar_demux_001_src24_data),          //           .data
		.src24_channel       (cmd_xbar_demux_001_src24_channel),       //           .channel
		.src24_startofpacket (cmd_xbar_demux_001_src24_startofpacket), //           .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_001_src24_endofpacket),   //           .endofpacket
		.src25_ready         (cmd_xbar_demux_001_src25_ready),         //      src25.ready
		.src25_valid         (cmd_xbar_demux_001_src25_valid),         //           .valid
		.src25_data          (cmd_xbar_demux_001_src25_data),          //           .data
		.src25_channel       (cmd_xbar_demux_001_src25_channel),       //           .channel
		.src25_startofpacket (cmd_xbar_demux_001_src25_startofpacket), //           .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_001_src25_endofpacket),   //           .endofpacket
		.src26_ready         (cmd_xbar_demux_001_src26_ready),         //      src26.ready
		.src26_valid         (cmd_xbar_demux_001_src26_valid),         //           .valid
		.src26_data          (cmd_xbar_demux_001_src26_data),          //           .data
		.src26_channel       (cmd_xbar_demux_001_src26_channel),       //           .channel
		.src26_startofpacket (cmd_xbar_demux_001_src26_startofpacket), //           .startofpacket
		.src26_endofpacket   (cmd_xbar_demux_001_src26_endofpacket),   //           .endofpacket
		.src27_ready         (cmd_xbar_demux_001_src27_ready),         //      src27.ready
		.src27_valid         (cmd_xbar_demux_001_src27_valid),         //           .valid
		.src27_data          (cmd_xbar_demux_001_src27_data),          //           .data
		.src27_channel       (cmd_xbar_demux_001_src27_channel),       //           .channel
		.src27_startofpacket (cmd_xbar_demux_001_src27_startofpacket), //           .startofpacket
		.src27_endofpacket   (cmd_xbar_demux_001_src27_endofpacket),   //           .endofpacket
		.src28_ready         (cmd_xbar_demux_001_src28_ready),         //      src28.ready
		.src28_valid         (cmd_xbar_demux_001_src28_valid),         //           .valid
		.src28_data          (cmd_xbar_demux_001_src28_data),          //           .data
		.src28_channel       (cmd_xbar_demux_001_src28_channel),       //           .channel
		.src28_startofpacket (cmd_xbar_demux_001_src28_startofpacket), //           .startofpacket
		.src28_endofpacket   (cmd_xbar_demux_001_src28_endofpacket),   //           .endofpacket
		.src29_ready         (cmd_xbar_demux_001_src29_ready),         //      src29.ready
		.src29_valid         (cmd_xbar_demux_001_src29_valid),         //           .valid
		.src29_data          (cmd_xbar_demux_001_src29_data),          //           .data
		.src29_channel       (cmd_xbar_demux_001_src29_channel),       //           .channel
		.src29_startofpacket (cmd_xbar_demux_001_src29_startofpacket), //           .startofpacket
		.src29_endofpacket   (cmd_xbar_demux_001_src29_endofpacket),   //           .endofpacket
		.src30_ready         (cmd_xbar_demux_001_src30_ready),         //      src30.ready
		.src30_valid         (cmd_xbar_demux_001_src30_valid),         //           .valid
		.src30_data          (cmd_xbar_demux_001_src30_data),          //           .data
		.src30_channel       (cmd_xbar_demux_001_src30_channel),       //           .channel
		.src30_startofpacket (cmd_xbar_demux_001_src30_startofpacket), //           .startofpacket
		.src30_endofpacket   (cmd_xbar_demux_001_src30_endofpacket),   //           .endofpacket
		.src31_ready         (cmd_xbar_demux_001_src31_ready),         //      src31.ready
		.src31_valid         (cmd_xbar_demux_001_src31_valid),         //           .valid
		.src31_data          (cmd_xbar_demux_001_src31_data),          //           .data
		.src31_channel       (cmd_xbar_demux_001_src31_channel),       //           .channel
		.src31_startofpacket (cmd_xbar_demux_001_src31_startofpacket), //           .startofpacket
		.src31_endofpacket   (cmd_xbar_demux_001_src31_endofpacket),   //           .endofpacket
		.src32_ready         (cmd_xbar_demux_001_src32_ready),         //      src32.ready
		.src32_valid         (cmd_xbar_demux_001_src32_valid),         //           .valid
		.src32_data          (cmd_xbar_demux_001_src32_data),          //           .data
		.src32_channel       (cmd_xbar_demux_001_src32_channel),       //           .channel
		.src32_startofpacket (cmd_xbar_demux_001_src32_startofpacket), //           .startofpacket
		.src32_endofpacket   (cmd_xbar_demux_001_src32_endofpacket),   //           .endofpacket
		.src33_ready         (cmd_xbar_demux_001_src33_ready),         //      src33.ready
		.src33_valid         (cmd_xbar_demux_001_src33_valid),         //           .valid
		.src33_data          (cmd_xbar_demux_001_src33_data),          //           .data
		.src33_channel       (cmd_xbar_demux_001_src33_channel),       //           .channel
		.src33_startofpacket (cmd_xbar_demux_001_src33_startofpacket), //           .startofpacket
		.src33_endofpacket   (cmd_xbar_demux_001_src33_endofpacket),   //           .endofpacket
		.src34_ready         (cmd_xbar_demux_001_src34_ready),         //      src34.ready
		.src34_valid         (cmd_xbar_demux_001_src34_valid),         //           .valid
		.src34_data          (cmd_xbar_demux_001_src34_data),          //           .data
		.src34_channel       (cmd_xbar_demux_001_src34_channel),       //           .channel
		.src34_startofpacket (cmd_xbar_demux_001_src34_startofpacket), //           .startofpacket
		.src34_endofpacket   (cmd_xbar_demux_001_src34_endofpacket),   //           .endofpacket
		.src35_ready         (cmd_xbar_demux_001_src35_ready),         //      src35.ready
		.src35_valid         (cmd_xbar_demux_001_src35_valid),         //           .valid
		.src35_data          (cmd_xbar_demux_001_src35_data),          //           .data
		.src35_channel       (cmd_xbar_demux_001_src35_channel),       //           .channel
		.src35_startofpacket (cmd_xbar_demux_001_src35_startofpacket), //           .startofpacket
		.src35_endofpacket   (cmd_xbar_demux_001_src35_endofpacket),   //           .endofpacket
		.src36_ready         (cmd_xbar_demux_001_src36_ready),         //      src36.ready
		.src36_valid         (cmd_xbar_demux_001_src36_valid),         //           .valid
		.src36_data          (cmd_xbar_demux_001_src36_data),          //           .data
		.src36_channel       (cmd_xbar_demux_001_src36_channel),       //           .channel
		.src36_startofpacket (cmd_xbar_demux_001_src36_startofpacket), //           .startofpacket
		.src36_endofpacket   (cmd_xbar_demux_001_src36_endofpacket)    //           .endofpacket
	);

	de2i_150_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux rsp_xbar_demux (
		.clk                (altpll_0_c0_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_011 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_012 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_013 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_014 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_015 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_016 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_017 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_018 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_019 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_020 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_021 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_022 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_023 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_024 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_025 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_026 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_027 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_028 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_029 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_030 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_031 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_031_src_ready),               //      sink.ready
		.sink_channel       (id_router_031_src_channel),             //          .channel
		.sink_data          (id_router_031_src_data),                //          .data
		.sink_startofpacket (id_router_031_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_031_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_031_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_032 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_032_src_ready),               //      sink.ready
		.sink_channel       (id_router_032_src_channel),             //          .channel
		.sink_data          (id_router_032_src_data),                //          .data
		.sink_startofpacket (id_router_032_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_032_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_032_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_033 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_033_src_ready),               //      sink.ready
		.sink_channel       (id_router_033_src_channel),             //          .channel
		.sink_data          (id_router_033_src_data),                //          .data
		.sink_startofpacket (id_router_033_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_033_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_033_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_033_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_033_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_034 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_034_src_ready),               //      sink.ready
		.sink_channel       (id_router_034_src_channel),             //          .channel
		.sink_data          (id_router_034_src_data),                //          .data
		.sink_startofpacket (id_router_034_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_034_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_034_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_034_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_034_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_035 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_035_src_ready),               //      sink.ready
		.sink_channel       (id_router_035_src_channel),             //          .channel
		.sink_data          (id_router_035_src_data),                //          .data
		.sink_startofpacket (id_router_035_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_035_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_035_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_035_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_035_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_demux_002 rsp_xbar_demux_036 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_036_src_ready),               //      sink.ready
		.sink_channel       (id_router_036_src_channel),             //          .channel
		.sink_data          (id_router_036_src_data),                //          .data
		.sink_startofpacket (id_router_036_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_036_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_036_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_036_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (altpll_0_c0_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	de2i_150_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (altpll_0_c0_clk),                       //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_023_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_024_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (crosser_002_out_ready),                 //    sink25.ready
		.sink25_valid         (crosser_002_out_valid),                 //          .valid
		.sink25_channel       (crosser_002_out_channel),               //          .channel
		.sink25_data          (crosser_002_out_data),                  //          .data
		.sink25_startofpacket (crosser_002_out_startofpacket),         //          .startofpacket
		.sink25_endofpacket   (crosser_002_out_endofpacket),           //          .endofpacket
		.sink26_ready         (rsp_xbar_demux_026_src0_ready),         //    sink26.ready
		.sink26_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink26_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink26_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.sink26_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink26_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink27_ready         (rsp_xbar_demux_027_src0_ready),         //    sink27.ready
		.sink27_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink27_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink27_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.sink27_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink27_endofpacket   (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink28_ready         (rsp_xbar_demux_028_src0_ready),         //    sink28.ready
		.sink28_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink28_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink28_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.sink28_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink28_endofpacket   (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.sink29_ready         (rsp_xbar_demux_029_src0_ready),         //    sink29.ready
		.sink29_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink29_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink29_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.sink29_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink29_endofpacket   (rsp_xbar_demux_029_src0_endofpacket),   //          .endofpacket
		.sink30_ready         (rsp_xbar_demux_030_src0_ready),         //    sink30.ready
		.sink30_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.sink30_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.sink30_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.sink30_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.sink30_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.sink31_ready         (rsp_xbar_demux_031_src0_ready),         //    sink31.ready
		.sink31_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.sink31_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.sink31_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.sink31_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.sink31_endofpacket   (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.sink32_ready         (crosser_003_out_ready),                 //    sink32.ready
		.sink32_valid         (crosser_003_out_valid),                 //          .valid
		.sink32_channel       (crosser_003_out_channel),               //          .channel
		.sink32_data          (crosser_003_out_data),                  //          .data
		.sink32_startofpacket (crosser_003_out_startofpacket),         //          .startofpacket
		.sink32_endofpacket   (crosser_003_out_endofpacket),           //          .endofpacket
		.sink33_ready         (rsp_xbar_demux_033_src0_ready),         //    sink33.ready
		.sink33_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.sink33_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.sink33_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.sink33_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.sink33_endofpacket   (rsp_xbar_demux_033_src0_endofpacket),   //          .endofpacket
		.sink34_ready         (rsp_xbar_demux_034_src0_ready),         //    sink34.ready
		.sink34_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.sink34_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.sink34_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.sink34_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.sink34_endofpacket   (rsp_xbar_demux_034_src0_endofpacket),   //          .endofpacket
		.sink35_ready         (rsp_xbar_demux_035_src0_ready),         //    sink35.ready
		.sink35_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.sink35_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.sink35_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.sink35_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.sink35_endofpacket   (rsp_xbar_demux_035_src0_endofpacket),   //          .endofpacket
		.sink36_ready         (rsp_xbar_demux_036_src0_ready),         //    sink36.ready
		.sink36_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.sink36_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.sink36_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.sink36_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.sink36_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (99),
		.BITS_PER_SYMBOL     (99),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (37),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_0_c0_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (clk_clk),                                //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src25_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src25_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src25_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src25_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src25_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src25_data),          //              .data
		.out_ready         (crosser_out_ready),                      //           out.ready
		.out_valid         (crosser_out_valid),                      //              .valid
		.out_startofpacket (crosser_out_startofpacket),              //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),                //              .endofpacket
		.out_channel       (crosser_out_channel),                    //              .channel
		.out_data          (crosser_out_data),                       //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (99),
		.BITS_PER_SYMBOL     (99),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (37),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (altpll_0_c0_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (clk_clk),                                //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src32_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src32_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src32_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src32_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src32_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src32_data),          //              .data
		.out_ready         (crosser_001_out_ready),                  //           out.ready
		.out_valid         (crosser_001_out_valid),                  //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_001_out_channel),                //              .channel
		.out_data          (crosser_001_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (99),
		.BITS_PER_SYMBOL     (99),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (37),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_025_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_025_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_025_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_025_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_025_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_025_src0_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (99),
		.BITS_PER_SYMBOL     (99),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (37),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_032_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_032_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_032_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_032_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_032_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_032_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	de2i_150_irq_mapper irq_mapper (
		.clk            (altpll_0_c0_clk),                //        clk.clk
		.reset          (rst_controller_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),       //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),       //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),       //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),       //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),       //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),       //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),       //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),       //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),       //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),       //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),      // receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq),      // receiver11.irq
		.receiver12_irq (irq_mapper_receiver12_irq),      // receiver12.irq
		.receiver13_irq (irq_mapper_receiver13_irq),      // receiver13.irq
		.receiver14_irq (irq_mapper_receiver14_irq),      // receiver14.irq
		.receiver15_irq (irq_mapper_receiver15_irq),      // receiver15.irq
		.receiver16_irq (irq_mapper_receiver16_irq),      // receiver16.irq
		.receiver17_irq (irq_mapper_receiver17_irq),      // receiver17.irq
		.receiver18_irq (irq_mapper_receiver18_irq),      // receiver18.irq
		.receiver19_irq (irq_mapper_receiver19_irq),      // receiver19.irq
		.receiver20_irq (irq_mapper_receiver20_irq),      // receiver20.irq
		.sender_irq     (nios2_qsys_d_irq_irq)            //     sender.irq
	);

endmodule
